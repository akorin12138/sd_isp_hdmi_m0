// Verilog netlist created by TD v5.0.30786
// Tue Mar 19 12:06:16 2024

`timescale 1ns / 1ps
module crc7_bram  // crc7_bram.v(14)
  (
  addra,
  clka,
  dia,
  wea,
  doa
  );

  input [7:0] addra;  // crc7_bram.v(29)
  input clka;  // crc7_bram.v(31)
  input [7:0] dia;  // crc7_bram.v(28)
  input wea;  // crc7_bram.v(30)
  output [7:0] doa;  // crc7_bram.v(26)

  parameter ADDR_WIDTH_A = 8;
  parameter ADDR_WIDTH_B = 8;
  parameter DATA_DEPTH_A = 256;
  parameter DATA_DEPTH_B = 256;
  parameter DATA_WIDTH_A = 8;
  parameter DATA_WIDTH_B = 8;
  parameter REGMODE_A = "NOREG";
  parameter WRITEMODE_A = "NORMAL";

  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=256;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h6E677C754A435851262F343D020B1019777E656C535A41483F362D241B120900),
    .INIT_01(256'h5C554E4778716A63141D060F3039222B454C575E6168737A0D041F1629203B32),
    .INIT_02(256'h0A0318112E273C35424B5059666F747D131A0108373E252C5B5249407F766D64),
    .INIT_03(256'h38312A231C150E077079626B545D464F2128333A050C171E69607B724D445F56),
    .INIT_04(256'h2F263D340B021910676E757C434A5158363F242D121B00097E776C655A534841),
    .INIT_05(256'h1D140F0639302B22555C474E7178636A040D161F2029323B4C455E5768617A73),
    .INIT_06(256'h4B4259506F667D74030A1118272E353C525B4049767F646D1A1308013E372C25),
    .INIT_07(256'h79706B625D544F463138232A151C070E6069727B444D565F28213A330C051E17),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_256x8_sub_000000_000 (
    .addra({2'b00,addra,3'b111}),
    .clka(clka),
    .dia({open_n69,dia}),
    .wea(wea),
    .doa({open_n84,doa}));

endmodule 

