module Reciprocal(
    input wire[7:0]     Average,    //均值
    output reg[31:0]    Recip       //倒数,1位整数位，31位小数位
);

    always @ (*)
        begin
            case(Average)
                8'd0: Recip = 32'b00000000000000000000000000000000;
                8'd1: Recip = 32'b10000000000000000000000000000000;
                8'd2: Recip = 32'b01000000000000000000000000000000;
                8'd3: Recip = 32'b00101010101010101010101010101010;
                8'd4: Recip = 32'b00100000000000000000000000000000;
                8'd5: Recip = 32'b00011001100110011001100110011001;
                8'd6: Recip = 32'b00010101010101010101010101010101;
                8'd7: Recip = 32'b00010010010010010010010010010010;
                8'd8: Recip = 32'b00010000000000000000000000000000;
                8'd9: Recip = 32'b00001110001110001110001110001110;
                8'd10: Recip = 32'b00001100110011001100110011001100;
                8'd11: Recip = 32'b00001011101000101110100010111010;
                8'd12: Recip = 32'b00001010101010101010101010101010;
                8'd13: Recip = 32'b00001001110110001001110110001001;
                8'd14: Recip = 32'b00001001001001001001001001001001;
                8'd15: Recip = 32'b00001000100010001000100010001000;
                8'd16: Recip = 32'b00001000000000000000000000000000;
                8'd17: Recip = 32'b00000111100001111000011110000111;
                8'd18: Recip = 32'b00000111000111000111000111000111;
                8'd19: Recip = 32'b00000110101111001010000110101111;
                8'd20: Recip = 32'b00000110011001100110011001100110;
                8'd21: Recip = 32'b00000110000110000110000110000110;
                8'd22: Recip = 32'b00000101110100010111010001011101;
                8'd23: Recip = 32'b00000101100100001011001000010110;
                8'd24: Recip = 32'b00000101010101010101010101010101;
                8'd25: Recip = 32'b00000101000111101011100001010001;
                8'd26: Recip = 32'b00000100111011000100111011000100;
                8'd27: Recip = 32'b00000100101111011010000100101111;
                8'd28: Recip = 32'b00000100100100100100100100100100;
                8'd29: Recip = 32'b00000100011010011110111001011000;
                8'd30: Recip = 32'b00000100010001000100010001000100;
                8'd31: Recip = 32'b00000100001000010000100001000010;
                8'd32: Recip = 32'b00000100000000000000000000000000;
                8'd33: Recip = 32'b00000011111000001111100000111110;
                8'd34: Recip = 32'b00000011110000111100001111000011;
                8'd35: Recip = 32'b00000011101010000011101010000011;
                8'd36: Recip = 32'b00000011100011100011100011100011;
                8'd37: Recip = 32'b00000011011101011001111100100010;
                8'd38: Recip = 32'b00000011010111100101000011010111;
                8'd39: Recip = 32'b00000011010010000011010010000011;
                8'd40: Recip = 32'b00000011001100110011001100110011;
                8'd41: Recip = 32'b00000011000111110011100000110001;
                8'd42: Recip = 32'b00000011000011000011000011000011;
                8'd43: Recip = 32'b00000010111110100000101111101000;
                8'd44: Recip = 32'b00000010111010001011101000101110;
                8'd45: Recip = 32'b00000010110110000010110110000010;
                8'd46: Recip = 32'b00000010110010000101100100001011;
                8'd47: Recip = 32'b00000010101110010011000100000101;
                8'd48: Recip = 32'b00000010101010101010101010101010;
                8'd49: Recip = 32'b00000010100111001011110000010100;
                8'd50: Recip = 32'b00000010100011110101110000101000;
                8'd51: Recip = 32'b00000010100000101000001010000010;
                8'd52: Recip = 32'b00000010011101100010011101100010;
                8'd53: Recip = 32'b00000010011010100100001110011111;
                8'd54: Recip = 32'b00000010010111101101000010010111;
                8'd55: Recip = 32'b00000010010100111100100000100101;
                8'd56: Recip = 32'b00000010010010010010010010010010;
                8'd57: Recip = 32'b00000010001111101110000010001111;
                8'd58: Recip = 32'b00000010001101001111011100101100;
                8'd59: Recip = 32'b00000010001010110110001111001011;
                8'd60: Recip = 32'b00000010001000100010001000100010;
                8'd61: Recip = 32'b00000010000110010010111000101001;
                8'd62: Recip = 32'b00000010000100001000010000100001;
                8'd63: Recip = 32'b00000010000010000010000010000010;
                8'd64: Recip = 32'b00000010000000000000000000000000;
                8'd65: Recip = 32'b00000001111110000001111110000001;
                8'd66: Recip = 32'b00000001111100000111110000011111;
                8'd67: Recip = 32'b00000001111010010001001100011010;
                8'd68: Recip = 32'b00000001111000011110000111100001;
                8'd69: Recip = 32'b00000001110110101110011000000111;
                8'd70: Recip = 32'b00000001110101000001110101000001;
                8'd71: Recip = 32'b00000001110011011000010101101000;
                8'd72: Recip = 32'b00000001110001110001110001110001;
                8'd73: Recip = 32'b00000001110000001110000001110000;
                8'd74: Recip = 32'b00000001101110101100111110010001;
                8'd75: Recip = 32'b00000001101101001110100000011011;
                8'd76: Recip = 32'b00000001101011110010100001101011;
                8'd77: Recip = 32'b00000001101010011000111011110110;
                8'd78: Recip = 32'b00000001101001000001101001000001;
                8'd79: Recip = 32'b00000001100111101100100011101001;
                8'd80: Recip = 32'b00000001100110011001100110011001;
                8'd81: Recip = 32'b00000001100101001000101100001111;
                8'd82: Recip = 32'b00000001100011111001110000011000;
                8'd83: Recip = 32'b00000001100010101100101110010000;
                8'd84: Recip = 32'b00000001100001100001100001100001;
                8'd85: Recip = 32'b00000001100000011000000110000001;
                8'd86: Recip = 32'b00000001011111010000010111110100;
                8'd87: Recip = 32'b00000001011110001010010011001000;
                8'd88: Recip = 32'b00000001011101000101110100010111;
                8'd89: Recip = 32'b00000001011100000010111000000101;
                8'd90: Recip = 32'b00000001011011000001011011000001;
                8'd91: Recip = 32'b00000001011010000001011010000001;
                8'd92: Recip = 32'b00000001011001000010110010000101;
                8'd93: Recip = 32'b00000001011000000101100000010110;
                8'd94: Recip = 32'b00000001010111001001100010000010;
                8'd95: Recip = 32'b00000001010110001110110100100011;
                8'd96: Recip = 32'b00000001010101010101010101010101;
                8'd97: Recip = 32'b00000001010100011101000001111110;
                8'd98: Recip = 32'b00000001010011100101111000001010;
                8'd99: Recip = 32'b00000001010010101111110101101010;
                8'd100: Recip = 32'b00000001010001111010111000010100;
                8'd101: Recip = 32'b00000001010001000110111110000110;
                8'd102: Recip = 32'b00000001010000010100000101000001;
                8'd103: Recip = 32'b00000001001111100010001011001011;
                8'd104: Recip = 32'b00000001001110110001001110110001;
                8'd105: Recip = 32'b00000001001110000001001110000001;
                8'd106: Recip = 32'b00000001001101010010000111001111;
                8'd107: Recip = 32'b00000001001100100011111000110100;
                8'd108: Recip = 32'b00000001001011110110100001001011;
                8'd109: Recip = 32'b00000001001011001001111110110100;
                8'd110: Recip = 32'b00000001001010011110010000010010;
                8'd111: Recip = 32'b00000001001001110011010100001011;
                8'd112: Recip = 32'b00000001001001001001001001001001;
                8'd113: Recip = 32'b00000001001000011111101101111000;
                8'd114: Recip = 32'b00000001000111110111000001000111;
                8'd115: Recip = 32'b00000001000111001111000001101010;
                8'd116: Recip = 32'b00000001000110100111101110010110;
                8'd117: Recip = 32'b00000001000110000001000110000001;
                8'd118: Recip = 32'b00000001000101011011000111100101;
                8'd119: Recip = 32'b00000001000100110101110010000001;
                8'd120: Recip = 32'b00000001000100010001000100010001;
                8'd121: Recip = 32'b00000001000011101100111101010110;
                8'd122: Recip = 32'b00000001000011001001011100010100;
                8'd123: Recip = 32'b00000001000010100110100000010000;
                8'd124: Recip = 32'b00000001000010000100001000010000;
                8'd125: Recip = 32'b00000001000001100010010011011101;
                8'd126: Recip = 32'b00000001000001000001000001000001;
                8'd127: Recip = 32'b00000001000000100000010000001000;
                8'd128: Recip = 32'b00000001000000000000000000000000;
                8'd129: Recip = 32'b00000000111111100000001111111000;
                8'd130: Recip = 32'b00000000111111000000111111000000;
                8'd131: Recip = 32'b00000000111110100010001100101100;
                8'd132: Recip = 32'b00000000111110000011111000001111;
                8'd133: Recip = 32'b00000000111101100110000000111101;
                8'd134: Recip = 32'b00000000111101001000100110001101;
                8'd135: Recip = 32'b00000000111100101011100111010110;
                8'd136: Recip = 32'b00000000111100001111000011110000;
                8'd137: Recip = 32'b00000000111011110010111010110111;
                8'd138: Recip = 32'b00000000111011010111001100000011;
                8'd139: Recip = 32'b00000000111010111011110110110010;
                8'd140: Recip = 32'b00000000111010100000111010100000;
                8'd141: Recip = 32'b00000000111010000110010110101100;
                8'd142: Recip = 32'b00000000111001101100001010110100;
                8'd143: Recip = 32'b00000000111001010010010110011000;
                8'd144: Recip = 32'b00000000111000111000111000111000;
                8'd145: Recip = 32'b00000000111000011111110001111000;
                8'd146: Recip = 32'b00000000111000000111000000111000;
                8'd147: Recip = 32'b00000000110111101110100101011100;
                8'd148: Recip = 32'b00000000110111010110011111001000;
                8'd149: Recip = 32'b00000000110110111110101101100001;
                8'd150: Recip = 32'b00000000110110100111010000001101;
                8'd151: Recip = 32'b00000000110110010000000110110010;
                8'd152: Recip = 32'b00000000110101111001010000110101;
                8'd153: Recip = 32'b00000000110101100010101110000000;
                8'd154: Recip = 32'b00000000110101001100011101111011;
                8'd155: Recip = 32'b00000000110100110110100000001101;
                8'd156: Recip = 32'b00000000110100100000110100100000;
                8'd157: Recip = 32'b00000000110100001011011010011111;
                8'd158: Recip = 32'b00000000110011110110010001110100;
                8'd159: Recip = 32'b00000000110011100001011010001010;
                8'd160: Recip = 32'b00000000110011001100110011001100;
                8'd161: Recip = 32'b00000000110010111000011100100111;
                8'd162: Recip = 32'b00000000110010100100010110000111;
                8'd163: Recip = 32'b00000000110010010000011111011010;
                8'd164: Recip = 32'b00000000110001111100111000001100;
                8'd165: Recip = 32'b00000000110001101001100000001100;
                8'd166: Recip = 32'b00000000110001010110010111001000;
                8'd167: Recip = 32'b00000000110001000011011100101111;
                8'd168: Recip = 32'b00000000110000110000110000110000;
                8'd169: Recip = 32'b00000000110000011110010010111011;
                8'd170: Recip = 32'b00000000110000001100000011000000;
                8'd171: Recip = 32'b00000000101111111010000000101111;
                8'd172: Recip = 32'b00000000101111101000001011111010;
                8'd173: Recip = 32'b00000000101111010110100100010000;
                8'd174: Recip = 32'b00000000101111000101001001100100;
                8'd175: Recip = 32'b00000000101110110011111011100111;
                8'd176: Recip = 32'b00000000101110100010111010001011;
                8'd177: Recip = 32'b00000000101110010010000101000011;
                8'd178: Recip = 32'b00000000101110000001011100000010;
                8'd179: Recip = 32'b00000000101101110000111110111011;
                8'd180: Recip = 32'b00000000101101100000101101100000;
                8'd181: Recip = 32'b00000000101101010000100111100110;
                8'd182: Recip = 32'b00000000101101000000101101000000;
                8'd183: Recip = 32'b00000000101100110000111101100011;
                8'd184: Recip = 32'b00000000101100100001011001000010;
                8'd185: Recip = 32'b00000000101100010001111111010011;
                8'd186: Recip = 32'b00000000101100000010110000001011;
                8'd187: Recip = 32'b00000000101011110011101011011101;
                8'd188: Recip = 32'b00000000101011100100110001000001;
                8'd189: Recip = 32'b00000000101011010110000000101011;
                8'd190: Recip = 32'b00000000101011000111011010010001;
                8'd191: Recip = 32'b00000000101010111000111101101001;
                8'd192: Recip = 32'b00000000101010101010101010101010;
                8'd193: Recip = 32'b00000000101010011100100001001010;
                8'd194: Recip = 32'b00000000101010001110100000111111;
                8'd195: Recip = 32'b00000000101010000000101010000000;
                8'd196: Recip = 32'b00000000101001110010111100000101;
                8'd197: Recip = 32'b00000000101001100101010111000100;
                8'd198: Recip = 32'b00000000101001010111111010110101;
                8'd199: Recip = 32'b00000000101001001010100111001111;
                8'd200: Recip = 32'b00000000101000111101011100001010;
                8'd201: Recip = 32'b00000000101000110000011001011110;
                8'd202: Recip = 32'b00000000101000100011011111000011;
                8'd203: Recip = 32'b00000000101000010110101100110001;
                8'd204: Recip = 32'b00000000101000001010000010100000;
                8'd205: Recip = 32'b00000000100111111101100000001001;
                8'd206: Recip = 32'b00000000100111110001000101100101;
                8'd207: Recip = 32'b00000000100111100100110010101101;
                8'd208: Recip = 32'b00000000100111011000100111011000;
                8'd209: Recip = 32'b00000000100111001100100011100001;
                8'd210: Recip = 32'b00000000100111000000100111000000;
                8'd211: Recip = 32'b00000000100110110100110001101111;
                8'd212: Recip = 32'b00000000100110101001000011100111;
                8'd213: Recip = 32'b00000000100110011101011100100010;
                8'd214: Recip = 32'b00000000100110010001111100011010;
                8'd215: Recip = 32'b00000000100110000110100011001000;
                8'd216: Recip = 32'b00000000100101111011010000100101;
                8'd217: Recip = 32'b00000000100101110000000100101110;
                8'd218: Recip = 32'b00000000100101100100111111011010;
                8'd219: Recip = 32'b00000000100101011010000000100101;
                8'd220: Recip = 32'b00000000100101001111001000001001;
                8'd221: Recip = 32'b00000000100101000100010110000000;
                8'd222: Recip = 32'b00000000100100111001101010000101;
                8'd223: Recip = 32'b00000000100100101111000100010011;
                8'd224: Recip = 32'b00000000100100100100100100100100;
                8'd225: Recip = 32'b00000000100100011010001010110011;
                8'd226: Recip = 32'b00000000100100001111110110111100;
                8'd227: Recip = 32'b00000000100100000101101000111000;
                8'd228: Recip = 32'b00000000100011111011100000100011;
                8'd229: Recip = 32'b00000000100011110001011101111001;
                8'd230: Recip = 32'b00000000100011100111100000110101;
                8'd231: Recip = 32'b00000000100011011101101001010010;
                8'd232: Recip = 32'b00000000100011010011110111001011;
                8'd233: Recip = 32'b00000000100011001010001010011100;
                8'd234: Recip = 32'b00000000100011000000100011000000;
                8'd235: Recip = 32'b00000000100010110111000000110100;
                8'd236: Recip = 32'b00000000100010101101100011110010;
                8'd237: Recip = 32'b00000000100010100100001011111000;
                8'd238: Recip = 32'b00000000100010011010111001000000;
                8'd239: Recip = 32'b00000000100010010001101011000111;
                8'd240: Recip = 32'b00000000100010001000100010001000;
                8'd241: Recip = 32'b00000000100001111111011110000000;
                8'd242: Recip = 32'b00000000100001110110011110101011;
                8'd243: Recip = 32'b00000000100001101101100100000101;
                8'd244: Recip = 32'b00000000100001100100101110001010;
                8'd245: Recip = 32'b00000000100001011011111100110111;
                8'd246: Recip = 32'b00000000100001010011010000001000;
                8'd247: Recip = 32'b00000000100001001010100111111001;
                8'd248: Recip = 32'b00000000100001000010000100001000;
                8'd249: Recip = 32'b00000000100000111001100100110000;
                8'd250: Recip = 32'b00000000100000110001001001101110;
                8'd251: Recip = 32'b00000000100000101000110010111111;
                8'd252: Recip = 32'b00000000100000100000100000100000;
                8'd253: Recip = 32'b00000000100000011000010010001101;
                8'd254: Recip = 32'b00000000100000010000001000000100;
                8'd255: Recip = 32'b00000000100000001000000010000000;
                default:Recip = 32'b00000000000000000000000000000000;
            endcase 
        end
endmodule