//12bits to 8bits
module log12bitsTo8bits
(
   input		[11:0]	Pre_Data,
   output	reg	[7:0]	Post_Data
);

always@(*)
begin
	case(Pre_Data)
	12'h00 : Post_Data = 8'h01; 
	12'h01 : Post_Data = 8'h02; 
	12'h02 : Post_Data = 8'h02; 
	12'h03 : Post_Data = 8'h03; 
	12'h04 : Post_Data = 8'h03; 
	12'h05 : Post_Data = 8'h03; 
	12'h06 : Post_Data = 8'h04; 
	12'h07 : Post_Data = 8'h04; 
	12'h08 : Post_Data = 8'h04; 
	12'h09 : Post_Data = 8'h05; 
	12'h0A : Post_Data = 8'h05; 
	12'h0B : Post_Data = 8'h05; 
	12'h0C : Post_Data = 8'h06; 
	12'h0D : Post_Data = 8'h06; 
	12'h0E : Post_Data = 8'h06; 
	12'h0F : Post_Data = 8'h06; 
	12'h10 : Post_Data = 8'h07; 
	12'h11 : Post_Data = 8'h07; 
	12'h12 : Post_Data = 8'h07; 
	12'h13 : Post_Data = 8'h07; 
	12'h14 : Post_Data = 8'h08; 
	12'h15 : Post_Data = 8'h08; 
	12'h16 : Post_Data = 8'h08; 
	12'h17 : Post_Data = 8'h08; 
	12'h18 : Post_Data = 8'h09; 
	12'h19 : Post_Data = 8'h09; 
	12'h1A : Post_Data = 8'h09; 
	12'h1B : Post_Data = 8'h09; 
	12'h1C : Post_Data = 8'h09; 
	12'h1D : Post_Data = 8'h0A; 
	12'h1E : Post_Data = 8'h0A; 
	12'h1F : Post_Data = 8'h0A; 
	12'h20 : Post_Data = 8'h0A; 
	12'h21 : Post_Data = 8'h0A; 
	12'h22 : Post_Data = 8'h0B; 
	12'h23 : Post_Data = 8'h0B; 
	12'h24 : Post_Data = 8'h0B; 
	12'h25 : Post_Data = 8'h0B; 
	12'h26 : Post_Data = 8'h0C; 
	12'h27 : Post_Data = 8'h0C; 
	12'h28 : Post_Data = 8'h0C; 
	12'h29 : Post_Data = 8'h0C; 
	12'h2A : Post_Data = 8'h0C; 
	12'h2B : Post_Data = 8'h0C; 
	12'h2C : Post_Data = 8'h0D; 
	12'h2D : Post_Data = 8'h0D; 
	12'h2E : Post_Data = 8'h0D; 
	12'h2F : Post_Data = 8'h0D; 
	12'h30 : Post_Data = 8'h0D; 
	12'h31 : Post_Data = 8'h0E; 
	12'h32 : Post_Data = 8'h0E; 
	12'h33 : Post_Data = 8'h0E; 
	12'h34 : Post_Data = 8'h0E; 
	12'h35 : Post_Data = 8'h0E; 
	12'h36 : Post_Data = 8'h0E; 
	12'h37 : Post_Data = 8'h0F; 
	12'h38 : Post_Data = 8'h0F; 
	12'h39 : Post_Data = 8'h0F; 
	12'h3A : Post_Data = 8'h0F; 
	12'h3B : Post_Data = 8'h0F; 
	12'h3C : Post_Data = 8'h0F; 
	12'h3D : Post_Data = 8'h10; 
	12'h3E : Post_Data = 8'h10; 
	12'h3F : Post_Data = 8'h10; 
	12'h40 : Post_Data = 8'h10; 
	12'h41 : Post_Data = 8'h10; 
	12'h42 : Post_Data = 8'h10; 
	12'h43 : Post_Data = 8'h11; 
	12'h44 : Post_Data = 8'h11; 
	12'h45 : Post_Data = 8'h11; 
	12'h46 : Post_Data = 8'h11; 
	12'h47 : Post_Data = 8'h11; 
	12'h48 : Post_Data = 8'h11; 
	12'h49 : Post_Data = 8'h12; 
	12'h4A : Post_Data = 8'h12; 
	12'h4B : Post_Data = 8'h12; 
	12'h4C : Post_Data = 8'h12; 
	12'h4D : Post_Data = 8'h12; 
	12'h4E : Post_Data = 8'h12; 
	12'h4F : Post_Data = 8'h13; 
	12'h50 : Post_Data = 8'h13; 
	12'h51 : Post_Data = 8'h13; 
	12'h52 : Post_Data = 8'h13; 
	12'h53 : Post_Data = 8'h13; 
	12'h54 : Post_Data = 8'h13; 
	12'h55 : Post_Data = 8'h13; 
	12'h56 : Post_Data = 8'h14; 
	12'h57 : Post_Data = 8'h14; 
	12'h58 : Post_Data = 8'h14; 
	12'h59 : Post_Data = 8'h14; 
	12'h5A : Post_Data = 8'h14; 
	12'h5B : Post_Data = 8'h14; 
	12'h5C : Post_Data = 8'h15; 
	12'h5D : Post_Data = 8'h15; 
	12'h5E : Post_Data = 8'h15; 
	12'h5F : Post_Data = 8'h15; 
	12'h60 : Post_Data = 8'h15; 
	12'h61 : Post_Data = 8'h15; 
	12'h62 : Post_Data = 8'h15; 
	12'h63 : Post_Data = 8'h16; 
	12'h64 : Post_Data = 8'h16; 
	12'h65 : Post_Data = 8'h16; 
	12'h66 : Post_Data = 8'h16; 
	12'h67 : Post_Data = 8'h16; 
	12'h68 : Post_Data = 8'h16; 
	12'h69 : Post_Data = 8'h16; 
	12'h6A : Post_Data = 8'h17; 
	12'h6B : Post_Data = 8'h17; 
	12'h6C : Post_Data = 8'h17; 
	12'h6D : Post_Data = 8'h17; 
	12'h6E : Post_Data = 8'h17; 
	12'h6F : Post_Data = 8'h17; 
	12'h70 : Post_Data = 8'h17; 
	12'h71 : Post_Data = 8'h18; 
	12'h72 : Post_Data = 8'h18; 
	12'h73 : Post_Data = 8'h18; 
	12'h74 : Post_Data = 8'h18; 
	12'h75 : Post_Data = 8'h18; 
	12'h76 : Post_Data = 8'h18; 
	12'h77 : Post_Data = 8'h18; 
	12'h78 : Post_Data = 8'h18; 
	12'h79 : Post_Data = 8'h19; 
	12'h7A : Post_Data = 8'h19; 
	12'h7B : Post_Data = 8'h19; 
	12'h7C : Post_Data = 8'h19; 
	12'h7D : Post_Data = 8'h19; 
	12'h7E : Post_Data = 8'h19; 
	12'h7F : Post_Data = 8'h19; 
	12'h80 : Post_Data = 8'h1A; 
	12'h81 : Post_Data = 8'h1A; 
	12'h82 : Post_Data = 8'h1A; 
	12'h83 : Post_Data = 8'h1A; 
	12'h84 : Post_Data = 8'h1A; 
	12'h85 : Post_Data = 8'h1A; 
	12'h86 : Post_Data = 8'h1A; 
	12'h87 : Post_Data = 8'h1A; 
	12'h88 : Post_Data = 8'h1B; 
	12'h89 : Post_Data = 8'h1B; 
	12'h8A : Post_Data = 8'h1B; 
	12'h8B : Post_Data = 8'h1B; 
	12'h8C : Post_Data = 8'h1B; 
	12'h8D : Post_Data = 8'h1B; 
	12'h8E : Post_Data = 8'h1B; 
	12'h8F : Post_Data = 8'h1B; 
	12'h90 : Post_Data = 8'h1C; 
	12'h91 : Post_Data = 8'h1C; 
	12'h92 : Post_Data = 8'h1C; 
	12'h93 : Post_Data = 8'h1C; 
	12'h94 : Post_Data = 8'h1C; 
	12'h95 : Post_Data = 8'h1C; 
	12'h96 : Post_Data = 8'h1C; 
	12'h97 : Post_Data = 8'h1C; 
	12'h98 : Post_Data = 8'h1D; 
	12'h99 : Post_Data = 8'h1D; 
	12'h9A : Post_Data = 8'h1D; 
	12'h9B : Post_Data = 8'h1D; 
	12'h9C : Post_Data = 8'h1D; 
	12'h9D : Post_Data = 8'h1D; 
	12'h9E : Post_Data = 8'h1D; 
	12'h9F : Post_Data = 8'h1D; 
	12'hA0 : Post_Data = 8'h1E; 
	12'hA1 : Post_Data = 8'h1E; 
	12'hA2 : Post_Data = 8'h1E; 
	12'hA3 : Post_Data = 8'h1E; 
	12'hA4 : Post_Data = 8'h1E; 
	12'hA5 : Post_Data = 8'h1E; 
	12'hA6 : Post_Data = 8'h1E; 
	12'hA7 : Post_Data = 8'h1E; 
	12'hA8 : Post_Data = 8'h1F; 
	12'hA9 : Post_Data = 8'h1F; 
	12'hAA : Post_Data = 8'h1F; 
	12'hAB : Post_Data = 8'h1F; 
	12'hAC : Post_Data = 8'h1F; 
	12'hAD : Post_Data = 8'h1F; 
	12'hAE : Post_Data = 8'h1F; 
	12'hAF : Post_Data = 8'h1F; 
	12'hB0 : Post_Data = 8'h20; 
	12'hB1 : Post_Data = 8'h20; 
	12'hB2 : Post_Data = 8'h20; 
	12'hB3 : Post_Data = 8'h20; 
	12'hB4 : Post_Data = 8'h20; 
	12'hB5 : Post_Data = 8'h20; 
	12'hB6 : Post_Data = 8'h20; 
	12'hB7 : Post_Data = 8'h20; 
	12'hB8 : Post_Data = 8'h20; 
	12'hB9 : Post_Data = 8'h21; 
	12'hBA : Post_Data = 8'h21; 
	12'hBB : Post_Data = 8'h21; 
	12'hBC : Post_Data = 8'h21; 
	12'hBD : Post_Data = 8'h21; 
	12'hBE : Post_Data = 8'h21; 
	12'hBF : Post_Data = 8'h21; 
	12'hC0 : Post_Data = 8'h21; 
	12'hC1 : Post_Data = 8'h22; 
	12'hC2 : Post_Data = 8'h22; 
	12'hC3 : Post_Data = 8'h22; 
	12'hC4 : Post_Data = 8'h22; 
	12'hC5 : Post_Data = 8'h22; 
	12'hC6 : Post_Data = 8'h22; 
	12'hC7 : Post_Data = 8'h22; 
	12'hC8 : Post_Data = 8'h22; 
	12'hC9 : Post_Data = 8'h22; 
	12'hCA : Post_Data = 8'h23; 
	12'hCB : Post_Data = 8'h23; 
	12'hCC : Post_Data = 8'h23; 
	12'hCD : Post_Data = 8'h23; 
	12'hCE : Post_Data = 8'h23; 
	12'hCF : Post_Data = 8'h23; 
	12'hD0 : Post_Data = 8'h23; 
	12'hD1 : Post_Data = 8'h23; 
	12'hD2 : Post_Data = 8'h23; 
	12'hD3 : Post_Data = 8'h24; 
	12'hD4 : Post_Data = 8'h24; 
	12'hD5 : Post_Data = 8'h24; 
	12'hD6 : Post_Data = 8'h24; 
	12'hD7 : Post_Data = 8'h24; 
	12'hD8 : Post_Data = 8'h24; 
	12'hD9 : Post_Data = 8'h24; 
	12'hDA : Post_Data = 8'h24; 
	12'hDB : Post_Data = 8'h24; 
	12'hDC : Post_Data = 8'h25; 
	12'hDD : Post_Data = 8'h25; 
	12'hDE : Post_Data = 8'h25; 
	12'hDF : Post_Data = 8'h25; 
	12'hE0 : Post_Data = 8'h25; 
	12'hE1 : Post_Data = 8'h25; 
	12'hE2 : Post_Data = 8'h25; 
	12'hE3 : Post_Data = 8'h25; 
	12'hE4 : Post_Data = 8'h25; 
	12'hE5 : Post_Data = 8'h26; 
	12'hE6 : Post_Data = 8'h26; 
	12'hE7 : Post_Data = 8'h26; 
	12'hE8 : Post_Data = 8'h26; 
	12'hE9 : Post_Data = 8'h26; 
	12'hEA : Post_Data = 8'h26; 
	12'hEB : Post_Data = 8'h26; 
	12'hEC : Post_Data = 8'h26; 
	12'hED : Post_Data = 8'h26; 
	12'hEE : Post_Data = 8'h27; 
	12'hEF : Post_Data = 8'h27; 
	12'hF0 : Post_Data = 8'h27; 
	12'hF1 : Post_Data = 8'h27; 
	12'hF2 : Post_Data = 8'h27; 
	12'hF3 : Post_Data = 8'h27; 
	12'hF4 : Post_Data = 8'h27; 
	12'hF5 : Post_Data = 8'h27; 
	12'hF6 : Post_Data = 8'h27; 
	12'hF7 : Post_Data = 8'h27; 
	12'hF8 : Post_Data = 8'h28; 
	12'hF9 : Post_Data = 8'h28; 
	12'hFA : Post_Data = 8'h28; 
	12'hFB : Post_Data = 8'h28; 
	12'hFC : Post_Data = 8'h28; 
	12'hFD : Post_Data = 8'h28; 
	12'hFE : Post_Data = 8'h28; 
	12'hFF : Post_Data = 8'h28; 
	12'h100 : Post_Data = 8'h28; 
	12'h101 : Post_Data = 8'h29; 
	12'h102 : Post_Data = 8'h29; 
	12'h103 : Post_Data = 8'h29; 
	12'h104 : Post_Data = 8'h29; 
	12'h105 : Post_Data = 8'h29; 
	12'h106 : Post_Data = 8'h29; 
	12'h107 : Post_Data = 8'h29; 
	12'h108 : Post_Data = 8'h29; 
	12'h109 : Post_Data = 8'h29; 
	12'h10A : Post_Data = 8'h29; 
	12'h10B : Post_Data = 8'h2A; 
	12'h10C : Post_Data = 8'h2A; 
	12'h10D : Post_Data = 8'h2A; 
	12'h10E : Post_Data = 8'h2A; 
	12'h10F : Post_Data = 8'h2A; 
	12'h110 : Post_Data = 8'h2A; 
	12'h111 : Post_Data = 8'h2A; 
	12'h112 : Post_Data = 8'h2A; 
	12'h113 : Post_Data = 8'h2A; 
	12'h114 : Post_Data = 8'h2A; 
	12'h115 : Post_Data = 8'h2B; 
	12'h116 : Post_Data = 8'h2B; 
	12'h117 : Post_Data = 8'h2B; 
	12'h118 : Post_Data = 8'h2B; 
	12'h119 : Post_Data = 8'h2B; 
	12'h11A : Post_Data = 8'h2B; 
	12'h11B : Post_Data = 8'h2B; 
	12'h11C : Post_Data = 8'h2B; 
	12'h11D : Post_Data = 8'h2B; 
	12'h11E : Post_Data = 8'h2C; 
	12'h11F : Post_Data = 8'h2C; 
	12'h120 : Post_Data = 8'h2C; 
	12'h121 : Post_Data = 8'h2C; 
	12'h122 : Post_Data = 8'h2C; 
	12'h123 : Post_Data = 8'h2C; 
	12'h124 : Post_Data = 8'h2C; 
	12'h125 : Post_Data = 8'h2C; 
	12'h126 : Post_Data = 8'h2C; 
	12'h127 : Post_Data = 8'h2C; 
	12'h128 : Post_Data = 8'h2D; 
	12'h129 : Post_Data = 8'h2D; 
	12'h12A : Post_Data = 8'h2D; 
	12'h12B : Post_Data = 8'h2D; 
	12'h12C : Post_Data = 8'h2D; 
	12'h12D : Post_Data = 8'h2D; 
	12'h12E : Post_Data = 8'h2D; 
	12'h12F : Post_Data = 8'h2D; 
	12'h130 : Post_Data = 8'h2D; 
	12'h131 : Post_Data = 8'h2D; 
	12'h132 : Post_Data = 8'h2E; 
	12'h133 : Post_Data = 8'h2E; 
	12'h134 : Post_Data = 8'h2E; 
	12'h135 : Post_Data = 8'h2E; 
	12'h136 : Post_Data = 8'h2E; 
	12'h137 : Post_Data = 8'h2E; 
	12'h138 : Post_Data = 8'h2E; 
	12'h139 : Post_Data = 8'h2E; 
	12'h13A : Post_Data = 8'h2E; 
	12'h13B : Post_Data = 8'h2E; 
	12'h13C : Post_Data = 8'h2E; 
	12'h13D : Post_Data = 8'h2F; 
	12'h13E : Post_Data = 8'h2F; 
	12'h13F : Post_Data = 8'h2F; 
	12'h140 : Post_Data = 8'h2F; 
	12'h141 : Post_Data = 8'h2F; 
	12'h142 : Post_Data = 8'h2F; 
	12'h143 : Post_Data = 8'h2F; 
	12'h144 : Post_Data = 8'h2F; 
	12'h145 : Post_Data = 8'h2F; 
	12'h146 : Post_Data = 8'h2F; 
	12'h147 : Post_Data = 8'h30; 
	12'h148 : Post_Data = 8'h30; 
	12'h149 : Post_Data = 8'h30; 
	12'h14A : Post_Data = 8'h30; 
	12'h14B : Post_Data = 8'h30; 
	12'h14C : Post_Data = 8'h30; 
	12'h14D : Post_Data = 8'h30; 
	12'h14E : Post_Data = 8'h30; 
	12'h14F : Post_Data = 8'h30; 
	12'h150 : Post_Data = 8'h30; 
	12'h151 : Post_Data = 8'h31; 
	12'h152 : Post_Data = 8'h31; 
	12'h153 : Post_Data = 8'h31; 
	12'h154 : Post_Data = 8'h31; 
	12'h155 : Post_Data = 8'h31; 
	12'h156 : Post_Data = 8'h31; 
	12'h157 : Post_Data = 8'h31; 
	12'h158 : Post_Data = 8'h31; 
	12'h159 : Post_Data = 8'h31; 
	12'h15A : Post_Data = 8'h31; 
	12'h15B : Post_Data = 8'h31; 
	12'h15C : Post_Data = 8'h32; 
	12'h15D : Post_Data = 8'h32; 
	12'h15E : Post_Data = 8'h32; 
	12'h15F : Post_Data = 8'h32; 
	12'h160 : Post_Data = 8'h32; 
	12'h161 : Post_Data = 8'h32; 
	12'h162 : Post_Data = 8'h32; 
	12'h163 : Post_Data = 8'h32; 
	12'h164 : Post_Data = 8'h32; 
	12'h165 : Post_Data = 8'h32; 
	12'h166 : Post_Data = 8'h33; 
	12'h167 : Post_Data = 8'h33; 
	12'h168 : Post_Data = 8'h33; 
	12'h169 : Post_Data = 8'h33; 
	12'h16A : Post_Data = 8'h33; 
	12'h16B : Post_Data = 8'h33; 
	12'h16C : Post_Data = 8'h33; 
	12'h16D : Post_Data = 8'h33; 
	12'h16E : Post_Data = 8'h33; 
	12'h16F : Post_Data = 8'h33; 
	12'h170 : Post_Data = 8'h33; 
	12'h171 : Post_Data = 8'h34; 
	12'h172 : Post_Data = 8'h34; 
	12'h173 : Post_Data = 8'h34; 
	12'h174 : Post_Data = 8'h34; 
	12'h175 : Post_Data = 8'h34; 
	12'h176 : Post_Data = 8'h34; 
	12'h177 : Post_Data = 8'h34; 
	12'h178 : Post_Data = 8'h34; 
	12'h179 : Post_Data = 8'h34; 
	12'h17A : Post_Data = 8'h34; 
	12'h17B : Post_Data = 8'h34; 
	12'h17C : Post_Data = 8'h35; 
	12'h17D : Post_Data = 8'h35; 
	12'h17E : Post_Data = 8'h35; 
	12'h17F : Post_Data = 8'h35; 
	12'h180 : Post_Data = 8'h35; 
	12'h181 : Post_Data = 8'h35; 
	12'h182 : Post_Data = 8'h35; 
	12'h183 : Post_Data = 8'h35; 
	12'h184 : Post_Data = 8'h35; 
	12'h185 : Post_Data = 8'h35; 
	12'h186 : Post_Data = 8'h35; 
	12'h187 : Post_Data = 8'h36; 
	12'h188 : Post_Data = 8'h36; 
	12'h189 : Post_Data = 8'h36; 
	12'h18A : Post_Data = 8'h36; 
	12'h18B : Post_Data = 8'h36; 
	12'h18C : Post_Data = 8'h36; 
	12'h18D : Post_Data = 8'h36; 
	12'h18E : Post_Data = 8'h36; 
	12'h18F : Post_Data = 8'h36; 
	12'h190 : Post_Data = 8'h36; 
	12'h191 : Post_Data = 8'h36; 
	12'h192 : Post_Data = 8'h37; 
	12'h193 : Post_Data = 8'h37; 
	12'h194 : Post_Data = 8'h37; 
	12'h195 : Post_Data = 8'h37; 
	12'h196 : Post_Data = 8'h37; 
	12'h197 : Post_Data = 8'h37; 
	12'h198 : Post_Data = 8'h37; 
	12'h199 : Post_Data = 8'h37; 
	12'h19A : Post_Data = 8'h37; 
	12'h19B : Post_Data = 8'h37; 
	12'h19C : Post_Data = 8'h37; 
	12'h19D : Post_Data = 8'h38; 
	12'h19E : Post_Data = 8'h38; 
	12'h19F : Post_Data = 8'h38; 
	12'h1A0 : Post_Data = 8'h38; 
	12'h1A1 : Post_Data = 8'h38; 
	12'h1A2 : Post_Data = 8'h38; 
	12'h1A3 : Post_Data = 8'h38; 
	12'h1A4 : Post_Data = 8'h38; 
	12'h1A5 : Post_Data = 8'h38; 
	12'h1A6 : Post_Data = 8'h38; 
	12'h1A7 : Post_Data = 8'h38; 
	12'h1A8 : Post_Data = 8'h39; 
	12'h1A9 : Post_Data = 8'h39; 
	12'h1AA : Post_Data = 8'h39; 
	12'h1AB : Post_Data = 8'h39; 
	12'h1AC : Post_Data = 8'h39; 
	12'h1AD : Post_Data = 8'h39; 
	12'h1AE : Post_Data = 8'h39; 
	12'h1AF : Post_Data = 8'h39; 
	12'h1B0 : Post_Data = 8'h39; 
	12'h1B1 : Post_Data = 8'h39; 
	12'h1B2 : Post_Data = 8'h39; 
	12'h1B3 : Post_Data = 8'h39; 
	12'h1B4 : Post_Data = 8'h3A; 
	12'h1B5 : Post_Data = 8'h3A; 
	12'h1B6 : Post_Data = 8'h3A; 
	12'h1B7 : Post_Data = 8'h3A; 
	12'h1B8 : Post_Data = 8'h3A; 
	12'h1B9 : Post_Data = 8'h3A; 
	12'h1BA : Post_Data = 8'h3A; 
	12'h1BB : Post_Data = 8'h3A; 
	12'h1BC : Post_Data = 8'h3A; 
	12'h1BD : Post_Data = 8'h3A; 
	12'h1BE : Post_Data = 8'h3A; 
	12'h1BF : Post_Data = 8'h3B; 
	12'h1C0 : Post_Data = 8'h3B; 
	12'h1C1 : Post_Data = 8'h3B; 
	12'h1C2 : Post_Data = 8'h3B; 
	12'h1C3 : Post_Data = 8'h3B; 
	12'h1C4 : Post_Data = 8'h3B; 
	12'h1C5 : Post_Data = 8'h3B; 
	12'h1C6 : Post_Data = 8'h3B; 
	12'h1C7 : Post_Data = 8'h3B; 
	12'h1C8 : Post_Data = 8'h3B; 
	12'h1C9 : Post_Data = 8'h3B; 
	12'h1CA : Post_Data = 8'h3C; 
	12'h1CB : Post_Data = 8'h3C; 
	12'h1CC : Post_Data = 8'h3C; 
	12'h1CD : Post_Data = 8'h3C; 
	12'h1CE : Post_Data = 8'h3C; 
	12'h1CF : Post_Data = 8'h3C; 
	12'h1D0 : Post_Data = 8'h3C; 
	12'h1D1 : Post_Data = 8'h3C; 
	12'h1D2 : Post_Data = 8'h3C; 
	12'h1D3 : Post_Data = 8'h3C; 
	12'h1D4 : Post_Data = 8'h3C; 
	12'h1D5 : Post_Data = 8'h3C; 
	12'h1D6 : Post_Data = 8'h3D; 
	12'h1D7 : Post_Data = 8'h3D; 
	12'h1D8 : Post_Data = 8'h3D; 
	12'h1D9 : Post_Data = 8'h3D; 
	12'h1DA : Post_Data = 8'h3D; 
	12'h1DB : Post_Data = 8'h3D; 
	12'h1DC : Post_Data = 8'h3D; 
	12'h1DD : Post_Data = 8'h3D; 
	12'h1DE : Post_Data = 8'h3D; 
	12'h1DF : Post_Data = 8'h3D; 
	12'h1E0 : Post_Data = 8'h3D; 
	12'h1E1 : Post_Data = 8'h3D; 
	12'h1E2 : Post_Data = 8'h3E; 
	12'h1E3 : Post_Data = 8'h3E; 
	12'h1E4 : Post_Data = 8'h3E; 
	12'h1E5 : Post_Data = 8'h3E; 
	12'h1E6 : Post_Data = 8'h3E; 
	12'h1E7 : Post_Data = 8'h3E; 
	12'h1E8 : Post_Data = 8'h3E; 
	12'h1E9 : Post_Data = 8'h3E; 
	12'h1EA : Post_Data = 8'h3E; 
	12'h1EB : Post_Data = 8'h3E; 
	12'h1EC : Post_Data = 8'h3E; 
	12'h1ED : Post_Data = 8'h3E; 
	12'h1EE : Post_Data = 8'h3F; 
	12'h1EF : Post_Data = 8'h3F; 
	12'h1F0 : Post_Data = 8'h3F; 
	12'h1F1 : Post_Data = 8'h3F; 
	12'h1F2 : Post_Data = 8'h3F; 
	12'h1F3 : Post_Data = 8'h3F; 
	12'h1F4 : Post_Data = 8'h3F; 
	12'h1F5 : Post_Data = 8'h3F; 
	12'h1F6 : Post_Data = 8'h3F; 
	12'h1F7 : Post_Data = 8'h3F; 
	12'h1F8 : Post_Data = 8'h3F; 
	12'h1F9 : Post_Data = 8'h3F; 
	12'h1FA : Post_Data = 8'h40; 
	12'h1FB : Post_Data = 8'h40; 
	12'h1FC : Post_Data = 8'h40; 
	12'h1FD : Post_Data = 8'h40; 
	12'h1FE : Post_Data = 8'h40; 
	12'h1FF : Post_Data = 8'h40; 
	12'h200 : Post_Data = 8'h40; 
	12'h201 : Post_Data = 8'h40; 
	12'h202 : Post_Data = 8'h40; 
	12'h203 : Post_Data = 8'h40; 
	12'h204 : Post_Data = 8'h40; 
	12'h205 : Post_Data = 8'h40; 
	12'h206 : Post_Data = 8'h41; 
	12'h207 : Post_Data = 8'h41; 
	12'h208 : Post_Data = 8'h41; 
	12'h209 : Post_Data = 8'h41; 
	12'h20A : Post_Data = 8'h41; 
	12'h20B : Post_Data = 8'h41; 
	12'h20C : Post_Data = 8'h41; 
	12'h20D : Post_Data = 8'h41; 
	12'h20E : Post_Data = 8'h41; 
	12'h20F : Post_Data = 8'h41; 
	12'h210 : Post_Data = 8'h41; 
	12'h211 : Post_Data = 8'h41; 
	12'h212 : Post_Data = 8'h42; 
	12'h213 : Post_Data = 8'h42; 
	12'h214 : Post_Data = 8'h42; 
	12'h215 : Post_Data = 8'h42; 
	12'h216 : Post_Data = 8'h42; 
	12'h217 : Post_Data = 8'h42; 
	12'h218 : Post_Data = 8'h42; 
	12'h219 : Post_Data = 8'h42; 
	12'h21A : Post_Data = 8'h42; 
	12'h21B : Post_Data = 8'h42; 
	12'h21C : Post_Data = 8'h42; 
	12'h21D : Post_Data = 8'h42; 
	12'h21E : Post_Data = 8'h43; 
	12'h21F : Post_Data = 8'h43; 
	12'h220 : Post_Data = 8'h43; 
	12'h221 : Post_Data = 8'h43; 
	12'h222 : Post_Data = 8'h43; 
	12'h223 : Post_Data = 8'h43; 
	12'h224 : Post_Data = 8'h43; 
	12'h225 : Post_Data = 8'h43; 
	12'h226 : Post_Data = 8'h43; 
	12'h227 : Post_Data = 8'h43; 
	12'h228 : Post_Data = 8'h43; 
	12'h229 : Post_Data = 8'h43; 
	12'h22A : Post_Data = 8'h44; 
	12'h22B : Post_Data = 8'h44; 
	12'h22C : Post_Data = 8'h44; 
	12'h22D : Post_Data = 8'h44; 
	12'h22E : Post_Data = 8'h44; 
	12'h22F : Post_Data = 8'h44; 
	12'h230 : Post_Data = 8'h44; 
	12'h231 : Post_Data = 8'h44; 
	12'h232 : Post_Data = 8'h44; 
	12'h233 : Post_Data = 8'h44; 
	12'h234 : Post_Data = 8'h44; 
	12'h235 : Post_Data = 8'h44; 
	12'h236 : Post_Data = 8'h45; 
	12'h237 : Post_Data = 8'h45; 
	12'h238 : Post_Data = 8'h45; 
	12'h239 : Post_Data = 8'h45; 
	12'h23A : Post_Data = 8'h45; 
	12'h23B : Post_Data = 8'h45; 
	12'h23C : Post_Data = 8'h45; 
	12'h23D : Post_Data = 8'h45; 
	12'h23E : Post_Data = 8'h45; 
	12'h23F : Post_Data = 8'h45; 
	12'h240 : Post_Data = 8'h45; 
	12'h241 : Post_Data = 8'h45; 
	12'h242 : Post_Data = 8'h45; 
	12'h243 : Post_Data = 8'h46; 
	12'h244 : Post_Data = 8'h46; 
	12'h245 : Post_Data = 8'h46; 
	12'h246 : Post_Data = 8'h46; 
	12'h247 : Post_Data = 8'h46; 
	12'h248 : Post_Data = 8'h46; 
	12'h249 : Post_Data = 8'h46; 
	12'h24A : Post_Data = 8'h46; 
	12'h24B : Post_Data = 8'h46; 
	12'h24C : Post_Data = 8'h46; 
	12'h24D : Post_Data = 8'h46; 
	12'h24E : Post_Data = 8'h46; 
	12'h24F : Post_Data = 8'h47; 
	12'h250 : Post_Data = 8'h47; 
	12'h251 : Post_Data = 8'h47; 
	12'h252 : Post_Data = 8'h47; 
	12'h253 : Post_Data = 8'h47; 
	12'h254 : Post_Data = 8'h47; 
	12'h255 : Post_Data = 8'h47; 
	12'h256 : Post_Data = 8'h47; 
	12'h257 : Post_Data = 8'h47; 
	12'h258 : Post_Data = 8'h47; 
	12'h259 : Post_Data = 8'h47; 
	12'h25A : Post_Data = 8'h47; 
	12'h25B : Post_Data = 8'h47; 
	12'h25C : Post_Data = 8'h48; 
	12'h25D : Post_Data = 8'h48; 
	12'h25E : Post_Data = 8'h48; 
	12'h25F : Post_Data = 8'h48; 
	12'h260 : Post_Data = 8'h48; 
	12'h261 : Post_Data = 8'h48; 
	12'h262 : Post_Data = 8'h48; 
	12'h263 : Post_Data = 8'h48; 
	12'h264 : Post_Data = 8'h48; 
	12'h265 : Post_Data = 8'h48; 
	12'h266 : Post_Data = 8'h48; 
	12'h267 : Post_Data = 8'h48; 
	12'h268 : Post_Data = 8'h48; 
	12'h269 : Post_Data = 8'h49; 
	12'h26A : Post_Data = 8'h49; 
	12'h26B : Post_Data = 8'h49; 
	12'h26C : Post_Data = 8'h49; 
	12'h26D : Post_Data = 8'h49; 
	12'h26E : Post_Data = 8'h49; 
	12'h26F : Post_Data = 8'h49; 
	12'h270 : Post_Data = 8'h49; 
	12'h271 : Post_Data = 8'h49; 
	12'h272 : Post_Data = 8'h49; 
	12'h273 : Post_Data = 8'h49; 
	12'h274 : Post_Data = 8'h49; 
	12'h275 : Post_Data = 8'h49; 
	12'h276 : Post_Data = 8'h4A; 
	12'h277 : Post_Data = 8'h4A; 
	12'h278 : Post_Data = 8'h4A; 
	12'h279 : Post_Data = 8'h4A; 
	12'h27A : Post_Data = 8'h4A; 
	12'h27B : Post_Data = 8'h4A; 
	12'h27C : Post_Data = 8'h4A; 
	12'h27D : Post_Data = 8'h4A; 
	12'h27E : Post_Data = 8'h4A; 
	12'h27F : Post_Data = 8'h4A; 
	12'h280 : Post_Data = 8'h4A; 
	12'h281 : Post_Data = 8'h4A; 
	12'h282 : Post_Data = 8'h4A; 
	12'h283 : Post_Data = 8'h4B; 
	12'h284 : Post_Data = 8'h4B; 
	12'h285 : Post_Data = 8'h4B; 
	12'h286 : Post_Data = 8'h4B; 
	12'h287 : Post_Data = 8'h4B; 
	12'h288 : Post_Data = 8'h4B; 
	12'h289 : Post_Data = 8'h4B; 
	12'h28A : Post_Data = 8'h4B; 
	12'h28B : Post_Data = 8'h4B; 
	12'h28C : Post_Data = 8'h4B; 
	12'h28D : Post_Data = 8'h4B; 
	12'h28E : Post_Data = 8'h4B; 
	12'h28F : Post_Data = 8'h4B; 
	12'h290 : Post_Data = 8'h4C; 
	12'h291 : Post_Data = 8'h4C; 
	12'h292 : Post_Data = 8'h4C; 
	12'h293 : Post_Data = 8'h4C; 
	12'h294 : Post_Data = 8'h4C; 
	12'h295 : Post_Data = 8'h4C; 
	12'h296 : Post_Data = 8'h4C; 
	12'h297 : Post_Data = 8'h4C; 
	12'h298 : Post_Data = 8'h4C; 
	12'h299 : Post_Data = 8'h4C; 
	12'h29A : Post_Data = 8'h4C; 
	12'h29B : Post_Data = 8'h4C; 
	12'h29C : Post_Data = 8'h4C; 
	12'h29D : Post_Data = 8'h4D; 
	12'h29E : Post_Data = 8'h4D; 
	12'h29F : Post_Data = 8'h4D; 
	12'h2A0 : Post_Data = 8'h4D; 
	12'h2A1 : Post_Data = 8'h4D; 
	12'h2A2 : Post_Data = 8'h4D; 
	12'h2A3 : Post_Data = 8'h4D; 
	12'h2A4 : Post_Data = 8'h4D; 
	12'h2A5 : Post_Data = 8'h4D; 
	12'h2A6 : Post_Data = 8'h4D; 
	12'h2A7 : Post_Data = 8'h4D; 
	12'h2A8 : Post_Data = 8'h4D; 
	12'h2A9 : Post_Data = 8'h4D; 
	12'h2AA : Post_Data = 8'h4E; 
	12'h2AB : Post_Data = 8'h4E; 
	12'h2AC : Post_Data = 8'h4E; 
	12'h2AD : Post_Data = 8'h4E; 
	12'h2AE : Post_Data = 8'h4E; 
	12'h2AF : Post_Data = 8'h4E; 
	12'h2B0 : Post_Data = 8'h4E; 
	12'h2B1 : Post_Data = 8'h4E; 
	12'h2B2 : Post_Data = 8'h4E; 
	12'h2B3 : Post_Data = 8'h4E; 
	12'h2B4 : Post_Data = 8'h4E; 
	12'h2B5 : Post_Data = 8'h4E; 
	12'h2B6 : Post_Data = 8'h4E; 
	12'h2B7 : Post_Data = 8'h4F; 
	12'h2B8 : Post_Data = 8'h4F; 
	12'h2B9 : Post_Data = 8'h4F; 
	12'h2BA : Post_Data = 8'h4F; 
	12'h2BB : Post_Data = 8'h4F; 
	12'h2BC : Post_Data = 8'h4F; 
	12'h2BD : Post_Data = 8'h4F; 
	12'h2BE : Post_Data = 8'h4F; 
	12'h2BF : Post_Data = 8'h4F; 
	12'h2C0 : Post_Data = 8'h4F; 
	12'h2C1 : Post_Data = 8'h4F; 
	12'h2C2 : Post_Data = 8'h4F; 
	12'h2C3 : Post_Data = 8'h4F; 
	12'h2C4 : Post_Data = 8'h50; 
	12'h2C5 : Post_Data = 8'h50; 
	12'h2C6 : Post_Data = 8'h50; 
	12'h2C7 : Post_Data = 8'h50; 
	12'h2C8 : Post_Data = 8'h50; 
	12'h2C9 : Post_Data = 8'h50; 
	12'h2CA : Post_Data = 8'h50; 
	12'h2CB : Post_Data = 8'h50; 
	12'h2CC : Post_Data = 8'h50; 
	12'h2CD : Post_Data = 8'h50; 
	12'h2CE : Post_Data = 8'h50; 
	12'h2CF : Post_Data = 8'h50; 
	12'h2D0 : Post_Data = 8'h50; 
	12'h2D1 : Post_Data = 8'h50; 
	12'h2D2 : Post_Data = 8'h51; 
	12'h2D3 : Post_Data = 8'h51; 
	12'h2D4 : Post_Data = 8'h51; 
	12'h2D5 : Post_Data = 8'h51; 
	12'h2D6 : Post_Data = 8'h51; 
	12'h2D7 : Post_Data = 8'h51; 
	12'h2D8 : Post_Data = 8'h51; 
	12'h2D9 : Post_Data = 8'h51; 
	12'h2DA : Post_Data = 8'h51; 
	12'h2DB : Post_Data = 8'h51; 
	12'h2DC : Post_Data = 8'h51; 
	12'h2DD : Post_Data = 8'h51; 
	12'h2DE : Post_Data = 8'h51; 
	12'h2DF : Post_Data = 8'h52; 
	12'h2E0 : Post_Data = 8'h52; 
	12'h2E1 : Post_Data = 8'h52; 
	12'h2E2 : Post_Data = 8'h52; 
	12'h2E3 : Post_Data = 8'h52; 
	12'h2E4 : Post_Data = 8'h52; 
	12'h2E5 : Post_Data = 8'h52; 
	12'h2E6 : Post_Data = 8'h52; 
	12'h2E7 : Post_Data = 8'h52; 
	12'h2E8 : Post_Data = 8'h52; 
	12'h2E9 : Post_Data = 8'h52; 
	12'h2EA : Post_Data = 8'h52; 
	12'h2EB : Post_Data = 8'h52; 
	12'h2EC : Post_Data = 8'h52; 
	12'h2ED : Post_Data = 8'h53; 
	12'h2EE : Post_Data = 8'h53; 
	12'h2EF : Post_Data = 8'h53; 
	12'h2F0 : Post_Data = 8'h53; 
	12'h2F1 : Post_Data = 8'h53; 
	12'h2F2 : Post_Data = 8'h53; 
	12'h2F3 : Post_Data = 8'h53; 
	12'h2F4 : Post_Data = 8'h53; 
	12'h2F5 : Post_Data = 8'h53; 
	12'h2F6 : Post_Data = 8'h53; 
	12'h2F7 : Post_Data = 8'h53; 
	12'h2F8 : Post_Data = 8'h53; 
	12'h2F9 : Post_Data = 8'h53; 
	12'h2FA : Post_Data = 8'h53; 
	12'h2FB : Post_Data = 8'h54; 
	12'h2FC : Post_Data = 8'h54; 
	12'h2FD : Post_Data = 8'h54; 
	12'h2FE : Post_Data = 8'h54; 
	12'h2FF : Post_Data = 8'h54; 
	12'h300 : Post_Data = 8'h54; 
	12'h301 : Post_Data = 8'h54; 
	12'h302 : Post_Data = 8'h54; 
	12'h303 : Post_Data = 8'h54; 
	12'h304 : Post_Data = 8'h54; 
	12'h305 : Post_Data = 8'h54; 
	12'h306 : Post_Data = 8'h54; 
	12'h307 : Post_Data = 8'h54; 
	12'h308 : Post_Data = 8'h55; 
	12'h309 : Post_Data = 8'h55; 
	12'h30A : Post_Data = 8'h55; 
	12'h30B : Post_Data = 8'h55; 
	12'h30C : Post_Data = 8'h55; 
	12'h30D : Post_Data = 8'h55; 
	12'h30E : Post_Data = 8'h55; 
	12'h30F : Post_Data = 8'h55; 
	12'h310 : Post_Data = 8'h55; 
	12'h311 : Post_Data = 8'h55; 
	12'h312 : Post_Data = 8'h55; 
	12'h313 : Post_Data = 8'h55; 
	12'h314 : Post_Data = 8'h55; 
	12'h315 : Post_Data = 8'h55; 
	12'h316 : Post_Data = 8'h56; 
	12'h317 : Post_Data = 8'h56; 
	12'h318 : Post_Data = 8'h56; 
	12'h319 : Post_Data = 8'h56; 
	12'h31A : Post_Data = 8'h56; 
	12'h31B : Post_Data = 8'h56; 
	12'h31C : Post_Data = 8'h56; 
	12'h31D : Post_Data = 8'h56; 
	12'h31E : Post_Data = 8'h56; 
	12'h31F : Post_Data = 8'h56; 
	12'h320 : Post_Data = 8'h56; 
	12'h321 : Post_Data = 8'h56; 
	12'h322 : Post_Data = 8'h56; 
	12'h323 : Post_Data = 8'h56; 
	12'h324 : Post_Data = 8'h57; 
	12'h325 : Post_Data = 8'h57; 
	12'h326 : Post_Data = 8'h57; 
	12'h327 : Post_Data = 8'h57; 
	12'h328 : Post_Data = 8'h57; 
	12'h329 : Post_Data = 8'h57; 
	12'h32A : Post_Data = 8'h57; 
	12'h32B : Post_Data = 8'h57; 
	12'h32C : Post_Data = 8'h57; 
	12'h32D : Post_Data = 8'h57; 
	12'h32E : Post_Data = 8'h57; 
	12'h32F : Post_Data = 8'h57; 
	12'h330 : Post_Data = 8'h57; 
	12'h331 : Post_Data = 8'h57; 
	12'h332 : Post_Data = 8'h58; 
	12'h333 : Post_Data = 8'h58; 
	12'h334 : Post_Data = 8'h58; 
	12'h335 : Post_Data = 8'h58; 
	12'h336 : Post_Data = 8'h58; 
	12'h337 : Post_Data = 8'h58; 
	12'h338 : Post_Data = 8'h58; 
	12'h339 : Post_Data = 8'h58; 
	12'h33A : Post_Data = 8'h58; 
	12'h33B : Post_Data = 8'h58; 
	12'h33C : Post_Data = 8'h58; 
	12'h33D : Post_Data = 8'h58; 
	12'h33E : Post_Data = 8'h58; 
	12'h33F : Post_Data = 8'h58; 
	12'h340 : Post_Data = 8'h59; 
	12'h341 : Post_Data = 8'h59; 
	12'h342 : Post_Data = 8'h59; 
	12'h343 : Post_Data = 8'h59; 
	12'h344 : Post_Data = 8'h59; 
	12'h345 : Post_Data = 8'h59; 
	12'h346 : Post_Data = 8'h59; 
	12'h347 : Post_Data = 8'h59; 
	12'h348 : Post_Data = 8'h59; 
	12'h349 : Post_Data = 8'h59; 
	12'h34A : Post_Data = 8'h59; 
	12'h34B : Post_Data = 8'h59; 
	12'h34C : Post_Data = 8'h59; 
	12'h34D : Post_Data = 8'h59; 
	12'h34E : Post_Data = 8'h5A; 
	12'h34F : Post_Data = 8'h5A; 
	12'h350 : Post_Data = 8'h5A; 
	12'h351 : Post_Data = 8'h5A; 
	12'h352 : Post_Data = 8'h5A; 
	12'h353 : Post_Data = 8'h5A; 
	12'h354 : Post_Data = 8'h5A; 
	12'h355 : Post_Data = 8'h5A; 
	12'h356 : Post_Data = 8'h5A; 
	12'h357 : Post_Data = 8'h5A; 
	12'h358 : Post_Data = 8'h5A; 
	12'h359 : Post_Data = 8'h5A; 
	12'h35A : Post_Data = 8'h5A; 
	12'h35B : Post_Data = 8'h5A; 
	12'h35C : Post_Data = 8'h5B; 
	12'h35D : Post_Data = 8'h5B; 
	12'h35E : Post_Data = 8'h5B; 
	12'h35F : Post_Data = 8'h5B; 
	12'h360 : Post_Data = 8'h5B; 
	12'h361 : Post_Data = 8'h5B; 
	12'h362 : Post_Data = 8'h5B; 
	12'h363 : Post_Data = 8'h5B; 
	12'h364 : Post_Data = 8'h5B; 
	12'h365 : Post_Data = 8'h5B; 
	12'h366 : Post_Data = 8'h5B; 
	12'h367 : Post_Data = 8'h5B; 
	12'h368 : Post_Data = 8'h5B; 
	12'h369 : Post_Data = 8'h5B; 
	12'h36A : Post_Data = 8'h5B; 
	12'h36B : Post_Data = 8'h5C; 
	12'h36C : Post_Data = 8'h5C; 
	12'h36D : Post_Data = 8'h5C; 
	12'h36E : Post_Data = 8'h5C; 
	12'h36F : Post_Data = 8'h5C; 
	12'h370 : Post_Data = 8'h5C; 
	12'h371 : Post_Data = 8'h5C; 
	12'h372 : Post_Data = 8'h5C; 
	12'h373 : Post_Data = 8'h5C; 
	12'h374 : Post_Data = 8'h5C; 
	12'h375 : Post_Data = 8'h5C; 
	12'h376 : Post_Data = 8'h5C; 
	12'h377 : Post_Data = 8'h5C; 
	12'h378 : Post_Data = 8'h5C; 
	12'h379 : Post_Data = 8'h5D; 
	12'h37A : Post_Data = 8'h5D; 
	12'h37B : Post_Data = 8'h5D; 
	12'h37C : Post_Data = 8'h5D; 
	12'h37D : Post_Data = 8'h5D; 
	12'h37E : Post_Data = 8'h5D; 
	12'h37F : Post_Data = 8'h5D; 
	12'h380 : Post_Data = 8'h5D; 
	12'h381 : Post_Data = 8'h5D; 
	12'h382 : Post_Data = 8'h5D; 
	12'h383 : Post_Data = 8'h5D; 
	12'h384 : Post_Data = 8'h5D; 
	12'h385 : Post_Data = 8'h5D; 
	12'h386 : Post_Data = 8'h5D; 
	12'h387 : Post_Data = 8'h5D; 
	12'h388 : Post_Data = 8'h5E; 
	12'h389 : Post_Data = 8'h5E; 
	12'h38A : Post_Data = 8'h5E; 
	12'h38B : Post_Data = 8'h5E; 
	12'h38C : Post_Data = 8'h5E; 
	12'h38D : Post_Data = 8'h5E; 
	12'h38E : Post_Data = 8'h5E; 
	12'h38F : Post_Data = 8'h5E; 
	12'h390 : Post_Data = 8'h5E; 
	12'h391 : Post_Data = 8'h5E; 
	12'h392 : Post_Data = 8'h5E; 
	12'h393 : Post_Data = 8'h5E; 
	12'h394 : Post_Data = 8'h5E; 
	12'h395 : Post_Data = 8'h5E; 
	12'h396 : Post_Data = 8'h5F; 
	12'h397 : Post_Data = 8'h5F; 
	12'h398 : Post_Data = 8'h5F; 
	12'h399 : Post_Data = 8'h5F; 
	12'h39A : Post_Data = 8'h5F; 
	12'h39B : Post_Data = 8'h5F; 
	12'h39C : Post_Data = 8'h5F; 
	12'h39D : Post_Data = 8'h5F; 
	12'h39E : Post_Data = 8'h5F; 
	12'h39F : Post_Data = 8'h5F; 
	12'h3A0 : Post_Data = 8'h5F; 
	12'h3A1 : Post_Data = 8'h5F; 
	12'h3A2 : Post_Data = 8'h5F; 
	12'h3A3 : Post_Data = 8'h5F; 
	12'h3A4 : Post_Data = 8'h5F; 
	12'h3A5 : Post_Data = 8'h60; 
	12'h3A6 : Post_Data = 8'h60; 
	12'h3A7 : Post_Data = 8'h60; 
	12'h3A8 : Post_Data = 8'h60; 
	12'h3A9 : Post_Data = 8'h60; 
	12'h3AA : Post_Data = 8'h60; 
	12'h3AB : Post_Data = 8'h60; 
	12'h3AC : Post_Data = 8'h60; 
	12'h3AD : Post_Data = 8'h60; 
	12'h3AE : Post_Data = 8'h60; 
	12'h3AF : Post_Data = 8'h60; 
	12'h3B0 : Post_Data = 8'h60; 
	12'h3B1 : Post_Data = 8'h60; 
	12'h3B2 : Post_Data = 8'h60; 
	12'h3B3 : Post_Data = 8'h61; 
	12'h3B4 : Post_Data = 8'h61; 
	12'h3B5 : Post_Data = 8'h61; 
	12'h3B6 : Post_Data = 8'h61; 
	12'h3B7 : Post_Data = 8'h61; 
	12'h3B8 : Post_Data = 8'h61; 
	12'h3B9 : Post_Data = 8'h61; 
	12'h3BA : Post_Data = 8'h61; 
	12'h3BB : Post_Data = 8'h61; 
	12'h3BC : Post_Data = 8'h61; 
	12'h3BD : Post_Data = 8'h61; 
	12'h3BE : Post_Data = 8'h61; 
	12'h3BF : Post_Data = 8'h61; 
	12'h3C0 : Post_Data = 8'h61; 
	12'h3C1 : Post_Data = 8'h61; 
	12'h3C2 : Post_Data = 8'h62; 
	12'h3C3 : Post_Data = 8'h62; 
	12'h3C4 : Post_Data = 8'h62; 
	12'h3C5 : Post_Data = 8'h62; 
	12'h3C6 : Post_Data = 8'h62; 
	12'h3C7 : Post_Data = 8'h62; 
	12'h3C8 : Post_Data = 8'h62; 
	12'h3C9 : Post_Data = 8'h62; 
	12'h3CA : Post_Data = 8'h62; 
	12'h3CB : Post_Data = 8'h62; 
	12'h3CC : Post_Data = 8'h62; 
	12'h3CD : Post_Data = 8'h62; 
	12'h3CE : Post_Data = 8'h62; 
	12'h3CF : Post_Data = 8'h62; 
	12'h3D0 : Post_Data = 8'h62; 
	12'h3D1 : Post_Data = 8'h63; 
	12'h3D2 : Post_Data = 8'h63; 
	12'h3D3 : Post_Data = 8'h63; 
	12'h3D4 : Post_Data = 8'h63; 
	12'h3D5 : Post_Data = 8'h63; 
	12'h3D6 : Post_Data = 8'h63; 
	12'h3D7 : Post_Data = 8'h63; 
	12'h3D8 : Post_Data = 8'h63; 
	12'h3D9 : Post_Data = 8'h63; 
	12'h3DA : Post_Data = 8'h63; 
	12'h3DB : Post_Data = 8'h63; 
	12'h3DC : Post_Data = 8'h63; 
	12'h3DD : Post_Data = 8'h63; 
	12'h3DE : Post_Data = 8'h63; 
	12'h3DF : Post_Data = 8'h63; 
	12'h3E0 : Post_Data = 8'h64; 
	12'h3E1 : Post_Data = 8'h64; 
	12'h3E2 : Post_Data = 8'h64; 
	12'h3E3 : Post_Data = 8'h64; 
	12'h3E4 : Post_Data = 8'h64; 
	12'h3E5 : Post_Data = 8'h64; 
	12'h3E6 : Post_Data = 8'h64; 
	12'h3E7 : Post_Data = 8'h64; 
	12'h3E8 : Post_Data = 8'h64; 
	12'h3E9 : Post_Data = 8'h64; 
	12'h3EA : Post_Data = 8'h64; 
	12'h3EB : Post_Data = 8'h64; 
	12'h3EC : Post_Data = 8'h64; 
	12'h3ED : Post_Data = 8'h64; 
	12'h3EE : Post_Data = 8'h64; 
	12'h3EF : Post_Data = 8'h65; 
	12'h3F0 : Post_Data = 8'h65; 
	12'h3F1 : Post_Data = 8'h65; 
	12'h3F2 : Post_Data = 8'h65; 
	12'h3F3 : Post_Data = 8'h65; 
	12'h3F4 : Post_Data = 8'h65; 
	12'h3F5 : Post_Data = 8'h65; 
	12'h3F6 : Post_Data = 8'h65; 
	12'h3F7 : Post_Data = 8'h65; 
	12'h3F8 : Post_Data = 8'h65; 
	12'h3F9 : Post_Data = 8'h65; 
	12'h3FA : Post_Data = 8'h65; 
	12'h3FB : Post_Data = 8'h65; 
	12'h3FC : Post_Data = 8'h65; 
	12'h3FD : Post_Data = 8'h65; 
	12'h3FE : Post_Data = 8'h66; 
	12'h3FF : Post_Data = 8'h66; 
	12'h400 : Post_Data = 8'h66; 
	12'h401 : Post_Data = 8'h66; 
	12'h402 : Post_Data = 8'h66; 
	12'h403 : Post_Data = 8'h66; 
	12'h404 : Post_Data = 8'h66; 
	12'h405 : Post_Data = 8'h66; 
	12'h406 : Post_Data = 8'h66; 
	12'h407 : Post_Data = 8'h66; 
	12'h408 : Post_Data = 8'h66; 
	12'h409 : Post_Data = 8'h66; 
	12'h40A : Post_Data = 8'h66; 
	12'h40B : Post_Data = 8'h66; 
	12'h40C : Post_Data = 8'h66; 
	12'h40D : Post_Data = 8'h67; 
	12'h40E : Post_Data = 8'h67; 
	12'h40F : Post_Data = 8'h67; 
	12'h410 : Post_Data = 8'h67; 
	12'h411 : Post_Data = 8'h67; 
	12'h412 : Post_Data = 8'h67; 
	12'h413 : Post_Data = 8'h67; 
	12'h414 : Post_Data = 8'h67; 
	12'h415 : Post_Data = 8'h67; 
	12'h416 : Post_Data = 8'h67; 
	12'h417 : Post_Data = 8'h67; 
	12'h418 : Post_Data = 8'h67; 
	12'h419 : Post_Data = 8'h67; 
	12'h41A : Post_Data = 8'h67; 
	12'h41B : Post_Data = 8'h67; 
	12'h41C : Post_Data = 8'h68; 
	12'h41D : Post_Data = 8'h68; 
	12'h41E : Post_Data = 8'h68; 
	12'h41F : Post_Data = 8'h68; 
	12'h420 : Post_Data = 8'h68; 
	12'h421 : Post_Data = 8'h68; 
	12'h422 : Post_Data = 8'h68; 
	12'h423 : Post_Data = 8'h68; 
	12'h424 : Post_Data = 8'h68; 
	12'h425 : Post_Data = 8'h68; 
	12'h426 : Post_Data = 8'h68; 
	12'h427 : Post_Data = 8'h68; 
	12'h428 : Post_Data = 8'h68; 
	12'h429 : Post_Data = 8'h68; 
	12'h42A : Post_Data = 8'h68; 
	12'h42B : Post_Data = 8'h68; 
	12'h42C : Post_Data = 8'h69; 
	12'h42D : Post_Data = 8'h69; 
	12'h42E : Post_Data = 8'h69; 
	12'h42F : Post_Data = 8'h69; 
	12'h430 : Post_Data = 8'h69; 
	12'h431 : Post_Data = 8'h69; 
	12'h432 : Post_Data = 8'h69; 
	12'h433 : Post_Data = 8'h69; 
	12'h434 : Post_Data = 8'h69; 
	12'h435 : Post_Data = 8'h69; 
	12'h436 : Post_Data = 8'h69; 
	12'h437 : Post_Data = 8'h69; 
	12'h438 : Post_Data = 8'h69; 
	12'h439 : Post_Data = 8'h69; 
	12'h43A : Post_Data = 8'h69; 
	12'h43B : Post_Data = 8'h6A; 
	12'h43C : Post_Data = 8'h6A; 
	12'h43D : Post_Data = 8'h6A; 
	12'h43E : Post_Data = 8'h6A; 
	12'h43F : Post_Data = 8'h6A; 
	12'h440 : Post_Data = 8'h6A; 
	12'h441 : Post_Data = 8'h6A; 
	12'h442 : Post_Data = 8'h6A; 
	12'h443 : Post_Data = 8'h6A; 
	12'h444 : Post_Data = 8'h6A; 
	12'h445 : Post_Data = 8'h6A; 
	12'h446 : Post_Data = 8'h6A; 
	12'h447 : Post_Data = 8'h6A; 
	12'h448 : Post_Data = 8'h6A; 
	12'h449 : Post_Data = 8'h6A; 
	12'h44A : Post_Data = 8'h6A; 
	12'h44B : Post_Data = 8'h6B; 
	12'h44C : Post_Data = 8'h6B; 
	12'h44D : Post_Data = 8'h6B; 
	12'h44E : Post_Data = 8'h6B; 
	12'h44F : Post_Data = 8'h6B; 
	12'h450 : Post_Data = 8'h6B; 
	12'h451 : Post_Data = 8'h6B; 
	12'h452 : Post_Data = 8'h6B; 
	12'h453 : Post_Data = 8'h6B; 
	12'h454 : Post_Data = 8'h6B; 
	12'h455 : Post_Data = 8'h6B; 
	12'h456 : Post_Data = 8'h6B; 
	12'h457 : Post_Data = 8'h6B; 
	12'h458 : Post_Data = 8'h6B; 
	12'h459 : Post_Data = 8'h6B; 
	12'h45A : Post_Data = 8'h6C; 
	12'h45B : Post_Data = 8'h6C; 
	12'h45C : Post_Data = 8'h6C; 
	12'h45D : Post_Data = 8'h6C; 
	12'h45E : Post_Data = 8'h6C; 
	12'h45F : Post_Data = 8'h6C; 
	12'h460 : Post_Data = 8'h6C; 
	12'h461 : Post_Data = 8'h6C; 
	12'h462 : Post_Data = 8'h6C; 
	12'h463 : Post_Data = 8'h6C; 
	12'h464 : Post_Data = 8'h6C; 
	12'h465 : Post_Data = 8'h6C; 
	12'h466 : Post_Data = 8'h6C; 
	12'h467 : Post_Data = 8'h6C; 
	12'h468 : Post_Data = 8'h6C; 
	12'h469 : Post_Data = 8'h6C; 
	12'h46A : Post_Data = 8'h6D; 
	12'h46B : Post_Data = 8'h6D; 
	12'h46C : Post_Data = 8'h6D; 
	12'h46D : Post_Data = 8'h6D; 
	12'h46E : Post_Data = 8'h6D; 
	12'h46F : Post_Data = 8'h6D; 
	12'h470 : Post_Data = 8'h6D; 
	12'h471 : Post_Data = 8'h6D; 
	12'h472 : Post_Data = 8'h6D; 
	12'h473 : Post_Data = 8'h6D; 
	12'h474 : Post_Data = 8'h6D; 
	12'h475 : Post_Data = 8'h6D; 
	12'h476 : Post_Data = 8'h6D; 
	12'h477 : Post_Data = 8'h6D; 
	12'h478 : Post_Data = 8'h6D; 
	12'h479 : Post_Data = 8'h6E; 
	12'h47A : Post_Data = 8'h6E; 
	12'h47B : Post_Data = 8'h6E; 
	12'h47C : Post_Data = 8'h6E; 
	12'h47D : Post_Data = 8'h6E; 
	12'h47E : Post_Data = 8'h6E; 
	12'h47F : Post_Data = 8'h6E; 
	12'h480 : Post_Data = 8'h6E; 
	12'h481 : Post_Data = 8'h6E; 
	12'h482 : Post_Data = 8'h6E; 
	12'h483 : Post_Data = 8'h6E; 
	12'h484 : Post_Data = 8'h6E; 
	12'h485 : Post_Data = 8'h6E; 
	12'h486 : Post_Data = 8'h6E; 
	12'h487 : Post_Data = 8'h6E; 
	12'h488 : Post_Data = 8'h6E; 
	12'h489 : Post_Data = 8'h6F; 
	12'h48A : Post_Data = 8'h6F; 
	12'h48B : Post_Data = 8'h6F; 
	12'h48C : Post_Data = 8'h6F; 
	12'h48D : Post_Data = 8'h6F; 
	12'h48E : Post_Data = 8'h6F; 
	12'h48F : Post_Data = 8'h6F; 
	12'h490 : Post_Data = 8'h6F; 
	12'h491 : Post_Data = 8'h6F; 
	12'h492 : Post_Data = 8'h6F; 
	12'h493 : Post_Data = 8'h6F; 
	12'h494 : Post_Data = 8'h6F; 
	12'h495 : Post_Data = 8'h6F; 
	12'h496 : Post_Data = 8'h6F; 
	12'h497 : Post_Data = 8'h6F; 
	12'h498 : Post_Data = 8'h6F; 
	12'h499 : Post_Data = 8'h70; 
	12'h49A : Post_Data = 8'h70; 
	12'h49B : Post_Data = 8'h70; 
	12'h49C : Post_Data = 8'h70; 
	12'h49D : Post_Data = 8'h70; 
	12'h49E : Post_Data = 8'h70; 
	12'h49F : Post_Data = 8'h70; 
	12'h4A0 : Post_Data = 8'h70; 
	12'h4A1 : Post_Data = 8'h70; 
	12'h4A2 : Post_Data = 8'h70; 
	12'h4A3 : Post_Data = 8'h70; 
	12'h4A4 : Post_Data = 8'h70; 
	12'h4A5 : Post_Data = 8'h70; 
	12'h4A6 : Post_Data = 8'h70; 
	12'h4A7 : Post_Data = 8'h70; 
	12'h4A8 : Post_Data = 8'h70; 
	12'h4A9 : Post_Data = 8'h71; 
	12'h4AA : Post_Data = 8'h71; 
	12'h4AB : Post_Data = 8'h71; 
	12'h4AC : Post_Data = 8'h71; 
	12'h4AD : Post_Data = 8'h71; 
	12'h4AE : Post_Data = 8'h71; 
	12'h4AF : Post_Data = 8'h71; 
	12'h4B0 : Post_Data = 8'h71; 
	12'h4B1 : Post_Data = 8'h71; 
	12'h4B2 : Post_Data = 8'h71; 
	12'h4B3 : Post_Data = 8'h71; 
	12'h4B4 : Post_Data = 8'h71; 
	12'h4B5 : Post_Data = 8'h71; 
	12'h4B6 : Post_Data = 8'h71; 
	12'h4B7 : Post_Data = 8'h71; 
	12'h4B8 : Post_Data = 8'h71; 
	12'h4B9 : Post_Data = 8'h72; 
	12'h4BA : Post_Data = 8'h72; 
	12'h4BB : Post_Data = 8'h72; 
	12'h4BC : Post_Data = 8'h72; 
	12'h4BD : Post_Data = 8'h72; 
	12'h4BE : Post_Data = 8'h72; 
	12'h4BF : Post_Data = 8'h72; 
	12'h4C0 : Post_Data = 8'h72; 
	12'h4C1 : Post_Data = 8'h72; 
	12'h4C2 : Post_Data = 8'h72; 
	12'h4C3 : Post_Data = 8'h72; 
	12'h4C4 : Post_Data = 8'h72; 
	12'h4C5 : Post_Data = 8'h72; 
	12'h4C6 : Post_Data = 8'h72; 
	12'h4C7 : Post_Data = 8'h72; 
	12'h4C8 : Post_Data = 8'h72; 
	12'h4C9 : Post_Data = 8'h73; 
	12'h4CA : Post_Data = 8'h73; 
	12'h4CB : Post_Data = 8'h73; 
	12'h4CC : Post_Data = 8'h73; 
	12'h4CD : Post_Data = 8'h73; 
	12'h4CE : Post_Data = 8'h73; 
	12'h4CF : Post_Data = 8'h73; 
	12'h4D0 : Post_Data = 8'h73; 
	12'h4D1 : Post_Data = 8'h73; 
	12'h4D2 : Post_Data = 8'h73; 
	12'h4D3 : Post_Data = 8'h73; 
	12'h4D4 : Post_Data = 8'h73; 
	12'h4D5 : Post_Data = 8'h73; 
	12'h4D6 : Post_Data = 8'h73; 
	12'h4D7 : Post_Data = 8'h73; 
	12'h4D8 : Post_Data = 8'h73; 
	12'h4D9 : Post_Data = 8'h74; 
	12'h4DA : Post_Data = 8'h74; 
	12'h4DB : Post_Data = 8'h74; 
	12'h4DC : Post_Data = 8'h74; 
	12'h4DD : Post_Data = 8'h74; 
	12'h4DE : Post_Data = 8'h74; 
	12'h4DF : Post_Data = 8'h74; 
	12'h4E0 : Post_Data = 8'h74; 
	12'h4E1 : Post_Data = 8'h74; 
	12'h4E2 : Post_Data = 8'h74; 
	12'h4E3 : Post_Data = 8'h74; 
	12'h4E4 : Post_Data = 8'h74; 
	12'h4E5 : Post_Data = 8'h74; 
	12'h4E6 : Post_Data = 8'h74; 
	12'h4E7 : Post_Data = 8'h74; 
	12'h4E8 : Post_Data = 8'h74; 
	12'h4E9 : Post_Data = 8'h75; 
	12'h4EA : Post_Data = 8'h75; 
	12'h4EB : Post_Data = 8'h75; 
	12'h4EC : Post_Data = 8'h75; 
	12'h4ED : Post_Data = 8'h75; 
	12'h4EE : Post_Data = 8'h75; 
	12'h4EF : Post_Data = 8'h75; 
	12'h4F0 : Post_Data = 8'h75; 
	12'h4F1 : Post_Data = 8'h75; 
	12'h4F2 : Post_Data = 8'h75; 
	12'h4F3 : Post_Data = 8'h75; 
	12'h4F4 : Post_Data = 8'h75; 
	12'h4F5 : Post_Data = 8'h75; 
	12'h4F6 : Post_Data = 8'h75; 
	12'h4F7 : Post_Data = 8'h75; 
	12'h4F8 : Post_Data = 8'h75; 
	12'h4F9 : Post_Data = 8'h76; 
	12'h4FA : Post_Data = 8'h76; 
	12'h4FB : Post_Data = 8'h76; 
	12'h4FC : Post_Data = 8'h76; 
	12'h4FD : Post_Data = 8'h76; 
	12'h4FE : Post_Data = 8'h76; 
	12'h4FF : Post_Data = 8'h76; 
	12'h500 : Post_Data = 8'h76; 
	12'h501 : Post_Data = 8'h76; 
	12'h502 : Post_Data = 8'h76; 
	12'h503 : Post_Data = 8'h76; 
	12'h504 : Post_Data = 8'h76; 
	12'h505 : Post_Data = 8'h76; 
	12'h506 : Post_Data = 8'h76; 
	12'h507 : Post_Data = 8'h76; 
	12'h508 : Post_Data = 8'h76; 
	12'h509 : Post_Data = 8'h77; 
	12'h50A : Post_Data = 8'h77; 
	12'h50B : Post_Data = 8'h77; 
	12'h50C : Post_Data = 8'h77; 
	12'h50D : Post_Data = 8'h77; 
	12'h50E : Post_Data = 8'h77; 
	12'h50F : Post_Data = 8'h77; 
	12'h510 : Post_Data = 8'h77; 
	12'h511 : Post_Data = 8'h77; 
	12'h512 : Post_Data = 8'h77; 
	12'h513 : Post_Data = 8'h77; 
	12'h514 : Post_Data = 8'h77; 
	12'h515 : Post_Data = 8'h77; 
	12'h516 : Post_Data = 8'h77; 
	12'h517 : Post_Data = 8'h77; 
	12'h518 : Post_Data = 8'h77; 
	12'h519 : Post_Data = 8'h77; 
	12'h51A : Post_Data = 8'h78; 
	12'h51B : Post_Data = 8'h78; 
	12'h51C : Post_Data = 8'h78; 
	12'h51D : Post_Data = 8'h78; 
	12'h51E : Post_Data = 8'h78; 
	12'h51F : Post_Data = 8'h78; 
	12'h520 : Post_Data = 8'h78; 
	12'h521 : Post_Data = 8'h78; 
	12'h522 : Post_Data = 8'h78; 
	12'h523 : Post_Data = 8'h78; 
	12'h524 : Post_Data = 8'h78; 
	12'h525 : Post_Data = 8'h78; 
	12'h526 : Post_Data = 8'h78; 
	12'h527 : Post_Data = 8'h78; 
	12'h528 : Post_Data = 8'h78; 
	12'h529 : Post_Data = 8'h78; 
	12'h52A : Post_Data = 8'h79; 
	12'h52B : Post_Data = 8'h79; 
	12'h52C : Post_Data = 8'h79; 
	12'h52D : Post_Data = 8'h79; 
	12'h52E : Post_Data = 8'h79; 
	12'h52F : Post_Data = 8'h79; 
	12'h530 : Post_Data = 8'h79; 
	12'h531 : Post_Data = 8'h79; 
	12'h532 : Post_Data = 8'h79; 
	12'h533 : Post_Data = 8'h79; 
	12'h534 : Post_Data = 8'h79; 
	12'h535 : Post_Data = 8'h79; 
	12'h536 : Post_Data = 8'h79; 
	12'h537 : Post_Data = 8'h79; 
	12'h538 : Post_Data = 8'h79; 
	12'h539 : Post_Data = 8'h79; 
	12'h53A : Post_Data = 8'h79; 
	12'h53B : Post_Data = 8'h7A; 
	12'h53C : Post_Data = 8'h7A; 
	12'h53D : Post_Data = 8'h7A; 
	12'h53E : Post_Data = 8'h7A; 
	12'h53F : Post_Data = 8'h7A; 
	12'h540 : Post_Data = 8'h7A; 
	12'h541 : Post_Data = 8'h7A; 
	12'h542 : Post_Data = 8'h7A; 
	12'h543 : Post_Data = 8'h7A; 
	12'h544 : Post_Data = 8'h7A; 
	12'h545 : Post_Data = 8'h7A; 
	12'h546 : Post_Data = 8'h7A; 
	12'h547 : Post_Data = 8'h7A; 
	12'h548 : Post_Data = 8'h7A; 
	12'h549 : Post_Data = 8'h7A; 
	12'h54A : Post_Data = 8'h7A; 
	12'h54B : Post_Data = 8'h7B; 
	12'h54C : Post_Data = 8'h7B; 
	12'h54D : Post_Data = 8'h7B; 
	12'h54E : Post_Data = 8'h7B; 
	12'h54F : Post_Data = 8'h7B; 
	12'h550 : Post_Data = 8'h7B; 
	12'h551 : Post_Data = 8'h7B; 
	12'h552 : Post_Data = 8'h7B; 
	12'h553 : Post_Data = 8'h7B; 
	12'h554 : Post_Data = 8'h7B; 
	12'h555 : Post_Data = 8'h7B; 
	12'h556 : Post_Data = 8'h7B; 
	12'h557 : Post_Data = 8'h7B; 
	12'h558 : Post_Data = 8'h7B; 
	12'h559 : Post_Data = 8'h7B; 
	12'h55A : Post_Data = 8'h7B; 
	12'h55B : Post_Data = 8'h7B; 
	12'h55C : Post_Data = 8'h7C; 
	12'h55D : Post_Data = 8'h7C; 
	12'h55E : Post_Data = 8'h7C; 
	12'h55F : Post_Data = 8'h7C; 
	12'h560 : Post_Data = 8'h7C; 
	12'h561 : Post_Data = 8'h7C; 
	12'h562 : Post_Data = 8'h7C; 
	12'h563 : Post_Data = 8'h7C; 
	12'h564 : Post_Data = 8'h7C; 
	12'h565 : Post_Data = 8'h7C; 
	12'h566 : Post_Data = 8'h7C; 
	12'h567 : Post_Data = 8'h7C; 
	12'h568 : Post_Data = 8'h7C; 
	12'h569 : Post_Data = 8'h7C; 
	12'h56A : Post_Data = 8'h7C; 
	12'h56B : Post_Data = 8'h7C; 
	12'h56C : Post_Data = 8'h7C; 
	12'h56D : Post_Data = 8'h7D; 
	12'h56E : Post_Data = 8'h7D; 
	12'h56F : Post_Data = 8'h7D; 
	12'h570 : Post_Data = 8'h7D; 
	12'h571 : Post_Data = 8'h7D; 
	12'h572 : Post_Data = 8'h7D; 
	12'h573 : Post_Data = 8'h7D; 
	12'h574 : Post_Data = 8'h7D; 
	12'h575 : Post_Data = 8'h7D; 
	12'h576 : Post_Data = 8'h7D; 
	12'h577 : Post_Data = 8'h7D; 
	12'h578 : Post_Data = 8'h7D; 
	12'h579 : Post_Data = 8'h7D; 
	12'h57A : Post_Data = 8'h7D; 
	12'h57B : Post_Data = 8'h7D; 
	12'h57C : Post_Data = 8'h7D; 
	12'h57D : Post_Data = 8'h7E; 
	12'h57E : Post_Data = 8'h7E; 
	12'h57F : Post_Data = 8'h7E; 
	12'h580 : Post_Data = 8'h7E; 
	12'h581 : Post_Data = 8'h7E; 
	12'h582 : Post_Data = 8'h7E; 
	12'h583 : Post_Data = 8'h7E; 
	12'h584 : Post_Data = 8'h7E; 
	12'h585 : Post_Data = 8'h7E; 
	12'h586 : Post_Data = 8'h7E; 
	12'h587 : Post_Data = 8'h7E; 
	12'h588 : Post_Data = 8'h7E; 
	12'h589 : Post_Data = 8'h7E; 
	12'h58A : Post_Data = 8'h7E; 
	12'h58B : Post_Data = 8'h7E; 
	12'h58C : Post_Data = 8'h7E; 
	12'h58D : Post_Data = 8'h7E; 
	12'h58E : Post_Data = 8'h7F; 
	12'h58F : Post_Data = 8'h7F; 
	12'h590 : Post_Data = 8'h7F; 
	12'h591 : Post_Data = 8'h7F; 
	12'h592 : Post_Data = 8'h7F; 
	12'h593 : Post_Data = 8'h7F; 
	12'h594 : Post_Data = 8'h7F; 
	12'h595 : Post_Data = 8'h7F; 
	12'h596 : Post_Data = 8'h7F; 
	12'h597 : Post_Data = 8'h7F; 
	12'h598 : Post_Data = 8'h7F; 
	12'h599 : Post_Data = 8'h7F; 
	12'h59A : Post_Data = 8'h7F; 
	12'h59B : Post_Data = 8'h7F; 
	12'h59C : Post_Data = 8'h7F; 
	12'h59D : Post_Data = 8'h7F; 
	12'h59E : Post_Data = 8'h7F; 
	12'h59F : Post_Data = 8'h80; 
	12'h5A0 : Post_Data = 8'h80; 
	12'h5A1 : Post_Data = 8'h80; 
	12'h5A2 : Post_Data = 8'h80; 
	12'h5A3 : Post_Data = 8'h80; 
	12'h5A4 : Post_Data = 8'h80; 
	12'h5A5 : Post_Data = 8'h80; 
	12'h5A6 : Post_Data = 8'h80; 
	12'h5A7 : Post_Data = 8'h80; 
	12'h5A8 : Post_Data = 8'h80; 
	12'h5A9 : Post_Data = 8'h80; 
	12'h5AA : Post_Data = 8'h80; 
	12'h5AB : Post_Data = 8'h80; 
	12'h5AC : Post_Data = 8'h80; 
	12'h5AD : Post_Data = 8'h80; 
	12'h5AE : Post_Data = 8'h80; 
	12'h5AF : Post_Data = 8'h80; 
	12'h5B0 : Post_Data = 8'h81; 
	12'h5B1 : Post_Data = 8'h81; 
	12'h5B2 : Post_Data = 8'h81; 
	12'h5B3 : Post_Data = 8'h81; 
	12'h5B4 : Post_Data = 8'h81; 
	12'h5B5 : Post_Data = 8'h81; 
	12'h5B6 : Post_Data = 8'h81; 
	12'h5B7 : Post_Data = 8'h81; 
	12'h5B8 : Post_Data = 8'h81; 
	12'h5B9 : Post_Data = 8'h81; 
	12'h5BA : Post_Data = 8'h81; 
	12'h5BB : Post_Data = 8'h81; 
	12'h5BC : Post_Data = 8'h81; 
	12'h5BD : Post_Data = 8'h81; 
	12'h5BE : Post_Data = 8'h81; 
	12'h5BF : Post_Data = 8'h81; 
	12'h5C0 : Post_Data = 8'h81; 
	12'h5C1 : Post_Data = 8'h82; 
	12'h5C2 : Post_Data = 8'h82; 
	12'h5C3 : Post_Data = 8'h82; 
	12'h5C4 : Post_Data = 8'h82; 
	12'h5C5 : Post_Data = 8'h82; 
	12'h5C6 : Post_Data = 8'h82; 
	12'h5C7 : Post_Data = 8'h82; 
	12'h5C8 : Post_Data = 8'h82; 
	12'h5C9 : Post_Data = 8'h82; 
	12'h5CA : Post_Data = 8'h82; 
	12'h5CB : Post_Data = 8'h82; 
	12'h5CC : Post_Data = 8'h82; 
	12'h5CD : Post_Data = 8'h82; 
	12'h5CE : Post_Data = 8'h82; 
	12'h5CF : Post_Data = 8'h82; 
	12'h5D0 : Post_Data = 8'h82; 
	12'h5D1 : Post_Data = 8'h82; 
	12'h5D2 : Post_Data = 8'h83; 
	12'h5D3 : Post_Data = 8'h83; 
	12'h5D4 : Post_Data = 8'h83; 
	12'h5D5 : Post_Data = 8'h83; 
	12'h5D6 : Post_Data = 8'h83; 
	12'h5D7 : Post_Data = 8'h83; 
	12'h5D8 : Post_Data = 8'h83; 
	12'h5D9 : Post_Data = 8'h83; 
	12'h5DA : Post_Data = 8'h83; 
	12'h5DB : Post_Data = 8'h83; 
	12'h5DC : Post_Data = 8'h83; 
	12'h5DD : Post_Data = 8'h83; 
	12'h5DE : Post_Data = 8'h83; 
	12'h5DF : Post_Data = 8'h83; 
	12'h5E0 : Post_Data = 8'h83; 
	12'h5E1 : Post_Data = 8'h83; 
	12'h5E2 : Post_Data = 8'h83; 
	12'h5E3 : Post_Data = 8'h84; 
	12'h5E4 : Post_Data = 8'h84; 
	12'h5E5 : Post_Data = 8'h84; 
	12'h5E6 : Post_Data = 8'h84; 
	12'h5E7 : Post_Data = 8'h84; 
	12'h5E8 : Post_Data = 8'h84; 
	12'h5E9 : Post_Data = 8'h84; 
	12'h5EA : Post_Data = 8'h84; 
	12'h5EB : Post_Data = 8'h84; 
	12'h5EC : Post_Data = 8'h84; 
	12'h5ED : Post_Data = 8'h84; 
	12'h5EE : Post_Data = 8'h84; 
	12'h5EF : Post_Data = 8'h84; 
	12'h5F0 : Post_Data = 8'h84; 
	12'h5F1 : Post_Data = 8'h84; 
	12'h5F2 : Post_Data = 8'h84; 
	12'h5F3 : Post_Data = 8'h84; 
	12'h5F4 : Post_Data = 8'h84; 
	12'h5F5 : Post_Data = 8'h85; 
	12'h5F6 : Post_Data = 8'h85; 
	12'h5F7 : Post_Data = 8'h85; 
	12'h5F8 : Post_Data = 8'h85; 
	12'h5F9 : Post_Data = 8'h85; 
	12'h5FA : Post_Data = 8'h85; 
	12'h5FB : Post_Data = 8'h85; 
	12'h5FC : Post_Data = 8'h85; 
	12'h5FD : Post_Data = 8'h85; 
	12'h5FE : Post_Data = 8'h85; 
	12'h5FF : Post_Data = 8'h85; 
	12'h600 : Post_Data = 8'h85; 
	12'h601 : Post_Data = 8'h85; 
	12'h602 : Post_Data = 8'h85; 
	12'h603 : Post_Data = 8'h85; 
	12'h604 : Post_Data = 8'h85; 
	12'h605 : Post_Data = 8'h85; 
	12'h606 : Post_Data = 8'h86; 
	12'h607 : Post_Data = 8'h86; 
	12'h608 : Post_Data = 8'h86; 
	12'h609 : Post_Data = 8'h86; 
	12'h60A : Post_Data = 8'h86; 
	12'h60B : Post_Data = 8'h86; 
	12'h60C : Post_Data = 8'h86; 
	12'h60D : Post_Data = 8'h86; 
	12'h60E : Post_Data = 8'h86; 
	12'h60F : Post_Data = 8'h86; 
	12'h610 : Post_Data = 8'h86; 
	12'h611 : Post_Data = 8'h86; 
	12'h612 : Post_Data = 8'h86; 
	12'h613 : Post_Data = 8'h86; 
	12'h614 : Post_Data = 8'h86; 
	12'h615 : Post_Data = 8'h86; 
	12'h616 : Post_Data = 8'h86; 
	12'h617 : Post_Data = 8'h87; 
	12'h618 : Post_Data = 8'h87; 
	12'h619 : Post_Data = 8'h87; 
	12'h61A : Post_Data = 8'h87; 
	12'h61B : Post_Data = 8'h87; 
	12'h61C : Post_Data = 8'h87; 
	12'h61D : Post_Data = 8'h87; 
	12'h61E : Post_Data = 8'h87; 
	12'h61F : Post_Data = 8'h87; 
	12'h620 : Post_Data = 8'h87; 
	12'h621 : Post_Data = 8'h87; 
	12'h622 : Post_Data = 8'h87; 
	12'h623 : Post_Data = 8'h87; 
	12'h624 : Post_Data = 8'h87; 
	12'h625 : Post_Data = 8'h87; 
	12'h626 : Post_Data = 8'h87; 
	12'h627 : Post_Data = 8'h87; 
	12'h628 : Post_Data = 8'h87; 
	12'h629 : Post_Data = 8'h88; 
	12'h62A : Post_Data = 8'h88; 
	12'h62B : Post_Data = 8'h88; 
	12'h62C : Post_Data = 8'h88; 
	12'h62D : Post_Data = 8'h88; 
	12'h62E : Post_Data = 8'h88; 
	12'h62F : Post_Data = 8'h88; 
	12'h630 : Post_Data = 8'h88; 
	12'h631 : Post_Data = 8'h88; 
	12'h632 : Post_Data = 8'h88; 
	12'h633 : Post_Data = 8'h88; 
	12'h634 : Post_Data = 8'h88; 
	12'h635 : Post_Data = 8'h88; 
	12'h636 : Post_Data = 8'h88; 
	12'h637 : Post_Data = 8'h88; 
	12'h638 : Post_Data = 8'h88; 
	12'h639 : Post_Data = 8'h88; 
	12'h63A : Post_Data = 8'h89; 
	12'h63B : Post_Data = 8'h89; 
	12'h63C : Post_Data = 8'h89; 
	12'h63D : Post_Data = 8'h89; 
	12'h63E : Post_Data = 8'h89; 
	12'h63F : Post_Data = 8'h89; 
	12'h640 : Post_Data = 8'h89; 
	12'h641 : Post_Data = 8'h89; 
	12'h642 : Post_Data = 8'h89; 
	12'h643 : Post_Data = 8'h89; 
	12'h644 : Post_Data = 8'h89; 
	12'h645 : Post_Data = 8'h89; 
	12'h646 : Post_Data = 8'h89; 
	12'h647 : Post_Data = 8'h89; 
	12'h648 : Post_Data = 8'h89; 
	12'h649 : Post_Data = 8'h89; 
	12'h64A : Post_Data = 8'h89; 
	12'h64B : Post_Data = 8'h89; 
	12'h64C : Post_Data = 8'h8A; 
	12'h64D : Post_Data = 8'h8A; 
	12'h64E : Post_Data = 8'h8A; 
	12'h64F : Post_Data = 8'h8A; 
	12'h650 : Post_Data = 8'h8A; 
	12'h651 : Post_Data = 8'h8A; 
	12'h652 : Post_Data = 8'h8A; 
	12'h653 : Post_Data = 8'h8A; 
	12'h654 : Post_Data = 8'h8A; 
	12'h655 : Post_Data = 8'h8A; 
	12'h656 : Post_Data = 8'h8A; 
	12'h657 : Post_Data = 8'h8A; 
	12'h658 : Post_Data = 8'h8A; 
	12'h659 : Post_Data = 8'h8A; 
	12'h65A : Post_Data = 8'h8A; 
	12'h65B : Post_Data = 8'h8A; 
	12'h65C : Post_Data = 8'h8A; 
	12'h65D : Post_Data = 8'h8B; 
	12'h65E : Post_Data = 8'h8B; 
	12'h65F : Post_Data = 8'h8B; 
	12'h660 : Post_Data = 8'h8B; 
	12'h661 : Post_Data = 8'h8B; 
	12'h662 : Post_Data = 8'h8B; 
	12'h663 : Post_Data = 8'h8B; 
	12'h664 : Post_Data = 8'h8B; 
	12'h665 : Post_Data = 8'h8B; 
	12'h666 : Post_Data = 8'h8B; 
	12'h667 : Post_Data = 8'h8B; 
	12'h668 : Post_Data = 8'h8B; 
	12'h669 : Post_Data = 8'h8B; 
	12'h66A : Post_Data = 8'h8B; 
	12'h66B : Post_Data = 8'h8B; 
	12'h66C : Post_Data = 8'h8B; 
	12'h66D : Post_Data = 8'h8B; 
	12'h66E : Post_Data = 8'h8B; 
	12'h66F : Post_Data = 8'h8C; 
	12'h670 : Post_Data = 8'h8C; 
	12'h671 : Post_Data = 8'h8C; 
	12'h672 : Post_Data = 8'h8C; 
	12'h673 : Post_Data = 8'h8C; 
	12'h674 : Post_Data = 8'h8C; 
	12'h675 : Post_Data = 8'h8C; 
	12'h676 : Post_Data = 8'h8C; 
	12'h677 : Post_Data = 8'h8C; 
	12'h678 : Post_Data = 8'h8C; 
	12'h679 : Post_Data = 8'h8C; 
	12'h67A : Post_Data = 8'h8C; 
	12'h67B : Post_Data = 8'h8C; 
	12'h67C : Post_Data = 8'h8C; 
	12'h67D : Post_Data = 8'h8C; 
	12'h67E : Post_Data = 8'h8C; 
	12'h67F : Post_Data = 8'h8C; 
	12'h680 : Post_Data = 8'h8C; 
	12'h681 : Post_Data = 8'h8D; 
	12'h682 : Post_Data = 8'h8D; 
	12'h683 : Post_Data = 8'h8D; 
	12'h684 : Post_Data = 8'h8D; 
	12'h685 : Post_Data = 8'h8D; 
	12'h686 : Post_Data = 8'h8D; 
	12'h687 : Post_Data = 8'h8D; 
	12'h688 : Post_Data = 8'h8D; 
	12'h689 : Post_Data = 8'h8D; 
	12'h68A : Post_Data = 8'h8D; 
	12'h68B : Post_Data = 8'h8D; 
	12'h68C : Post_Data = 8'h8D; 
	12'h68D : Post_Data = 8'h8D; 
	12'h68E : Post_Data = 8'h8D; 
	12'h68F : Post_Data = 8'h8D; 
	12'h690 : Post_Data = 8'h8D; 
	12'h691 : Post_Data = 8'h8D; 
	12'h692 : Post_Data = 8'h8D; 
	12'h693 : Post_Data = 8'h8E; 
	12'h694 : Post_Data = 8'h8E; 
	12'h695 : Post_Data = 8'h8E; 
	12'h696 : Post_Data = 8'h8E; 
	12'h697 : Post_Data = 8'h8E; 
	12'h698 : Post_Data = 8'h8E; 
	12'h699 : Post_Data = 8'h8E; 
	12'h69A : Post_Data = 8'h8E; 
	12'h69B : Post_Data = 8'h8E; 
	12'h69C : Post_Data = 8'h8E; 
	12'h69D : Post_Data = 8'h8E; 
	12'h69E : Post_Data = 8'h8E; 
	12'h69F : Post_Data = 8'h8E; 
	12'h6A0 : Post_Data = 8'h8E; 
	12'h6A1 : Post_Data = 8'h8E; 
	12'h6A2 : Post_Data = 8'h8E; 
	12'h6A3 : Post_Data = 8'h8E; 
	12'h6A4 : Post_Data = 8'h8E; 
	12'h6A5 : Post_Data = 8'h8F; 
	12'h6A6 : Post_Data = 8'h8F; 
	12'h6A7 : Post_Data = 8'h8F; 
	12'h6A8 : Post_Data = 8'h8F; 
	12'h6A9 : Post_Data = 8'h8F; 
	12'h6AA : Post_Data = 8'h8F; 
	12'h6AB : Post_Data = 8'h8F; 
	12'h6AC : Post_Data = 8'h8F; 
	12'h6AD : Post_Data = 8'h8F; 
	12'h6AE : Post_Data = 8'h8F; 
	12'h6AF : Post_Data = 8'h8F; 
	12'h6B0 : Post_Data = 8'h8F; 
	12'h6B1 : Post_Data = 8'h8F; 
	12'h6B2 : Post_Data = 8'h8F; 
	12'h6B3 : Post_Data = 8'h8F; 
	12'h6B4 : Post_Data = 8'h8F; 
	12'h6B5 : Post_Data = 8'h8F; 
	12'h6B6 : Post_Data = 8'h8F; 
	12'h6B7 : Post_Data = 8'h90; 
	12'h6B8 : Post_Data = 8'h90; 
	12'h6B9 : Post_Data = 8'h90; 
	12'h6BA : Post_Data = 8'h90; 
	12'h6BB : Post_Data = 8'h90; 
	12'h6BC : Post_Data = 8'h90; 
	12'h6BD : Post_Data = 8'h90; 
	12'h6BE : Post_Data = 8'h90; 
	12'h6BF : Post_Data = 8'h90; 
	12'h6C0 : Post_Data = 8'h90; 
	12'h6C1 : Post_Data = 8'h90; 
	12'h6C2 : Post_Data = 8'h90; 
	12'h6C3 : Post_Data = 8'h90; 
	12'h6C4 : Post_Data = 8'h90; 
	12'h6C5 : Post_Data = 8'h90; 
	12'h6C6 : Post_Data = 8'h90; 
	12'h6C7 : Post_Data = 8'h90; 
	12'h6C8 : Post_Data = 8'h90; 
	12'h6C9 : Post_Data = 8'h91; 
	12'h6CA : Post_Data = 8'h91; 
	12'h6CB : Post_Data = 8'h91; 
	12'h6CC : Post_Data = 8'h91; 
	12'h6CD : Post_Data = 8'h91; 
	12'h6CE : Post_Data = 8'h91; 
	12'h6CF : Post_Data = 8'h91; 
	12'h6D0 : Post_Data = 8'h91; 
	12'h6D1 : Post_Data = 8'h91; 
	12'h6D2 : Post_Data = 8'h91; 
	12'h6D3 : Post_Data = 8'h91; 
	12'h6D4 : Post_Data = 8'h91; 
	12'h6D5 : Post_Data = 8'h91; 
	12'h6D6 : Post_Data = 8'h91; 
	12'h6D7 : Post_Data = 8'h91; 
	12'h6D8 : Post_Data = 8'h91; 
	12'h6D9 : Post_Data = 8'h91; 
	12'h6DA : Post_Data = 8'h91; 
	12'h6DB : Post_Data = 8'h92; 
	12'h6DC : Post_Data = 8'h92; 
	12'h6DD : Post_Data = 8'h92; 
	12'h6DE : Post_Data = 8'h92; 
	12'h6DF : Post_Data = 8'h92; 
	12'h6E0 : Post_Data = 8'h92; 
	12'h6E1 : Post_Data = 8'h92; 
	12'h6E2 : Post_Data = 8'h92; 
	12'h6E3 : Post_Data = 8'h92; 
	12'h6E4 : Post_Data = 8'h92; 
	12'h6E5 : Post_Data = 8'h92; 
	12'h6E6 : Post_Data = 8'h92; 
	12'h6E7 : Post_Data = 8'h92; 
	12'h6E8 : Post_Data = 8'h92; 
	12'h6E9 : Post_Data = 8'h92; 
	12'h6EA : Post_Data = 8'h92; 
	12'h6EB : Post_Data = 8'h92; 
	12'h6EC : Post_Data = 8'h92; 
	12'h6ED : Post_Data = 8'h93; 
	12'h6EE : Post_Data = 8'h93; 
	12'h6EF : Post_Data = 8'h93; 
	12'h6F0 : Post_Data = 8'h93; 
	12'h6F1 : Post_Data = 8'h93; 
	12'h6F2 : Post_Data = 8'h93; 
	12'h6F3 : Post_Data = 8'h93; 
	12'h6F4 : Post_Data = 8'h93; 
	12'h6F5 : Post_Data = 8'h93; 
	12'h6F6 : Post_Data = 8'h93; 
	12'h6F7 : Post_Data = 8'h93; 
	12'h6F8 : Post_Data = 8'h93; 
	12'h6F9 : Post_Data = 8'h93; 
	12'h6FA : Post_Data = 8'h93; 
	12'h6FB : Post_Data = 8'h93; 
	12'h6FC : Post_Data = 8'h93; 
	12'h6FD : Post_Data = 8'h93; 
	12'h6FE : Post_Data = 8'h93; 
	12'h6FF : Post_Data = 8'h94; 
	12'h700 : Post_Data = 8'h94; 
	12'h701 : Post_Data = 8'h94; 
	12'h702 : Post_Data = 8'h94; 
	12'h703 : Post_Data = 8'h94; 
	12'h704 : Post_Data = 8'h94; 
	12'h705 : Post_Data = 8'h94; 
	12'h706 : Post_Data = 8'h94; 
	12'h707 : Post_Data = 8'h94; 
	12'h708 : Post_Data = 8'h94; 
	12'h709 : Post_Data = 8'h94; 
	12'h70A : Post_Data = 8'h94; 
	12'h70B : Post_Data = 8'h94; 
	12'h70C : Post_Data = 8'h94; 
	12'h70D : Post_Data = 8'h94; 
	12'h70E : Post_Data = 8'h94; 
	12'h70F : Post_Data = 8'h94; 
	12'h710 : Post_Data = 8'h94; 
	12'h711 : Post_Data = 8'h95; 
	12'h712 : Post_Data = 8'h95; 
	12'h713 : Post_Data = 8'h95; 
	12'h714 : Post_Data = 8'h95; 
	12'h715 : Post_Data = 8'h95; 
	12'h716 : Post_Data = 8'h95; 
	12'h717 : Post_Data = 8'h95; 
	12'h718 : Post_Data = 8'h95; 
	12'h719 : Post_Data = 8'h95; 
	12'h71A : Post_Data = 8'h95; 
	12'h71B : Post_Data = 8'h95; 
	12'h71C : Post_Data = 8'h95; 
	12'h71D : Post_Data = 8'h95; 
	12'h71E : Post_Data = 8'h95; 
	12'h71F : Post_Data = 8'h95; 
	12'h720 : Post_Data = 8'h95; 
	12'h721 : Post_Data = 8'h95; 
	12'h722 : Post_Data = 8'h95; 
	12'h723 : Post_Data = 8'h96; 
	12'h724 : Post_Data = 8'h96; 
	12'h725 : Post_Data = 8'h96; 
	12'h726 : Post_Data = 8'h96; 
	12'h727 : Post_Data = 8'h96; 
	12'h728 : Post_Data = 8'h96; 
	12'h729 : Post_Data = 8'h96; 
	12'h72A : Post_Data = 8'h96; 
	12'h72B : Post_Data = 8'h96; 
	12'h72C : Post_Data = 8'h96; 
	12'h72D : Post_Data = 8'h96; 
	12'h72E : Post_Data = 8'h96; 
	12'h72F : Post_Data = 8'h96; 
	12'h730 : Post_Data = 8'h96; 
	12'h731 : Post_Data = 8'h96; 
	12'h732 : Post_Data = 8'h96; 
	12'h733 : Post_Data = 8'h96; 
	12'h734 : Post_Data = 8'h96; 
	12'h735 : Post_Data = 8'h96; 
	12'h736 : Post_Data = 8'h97; 
	12'h737 : Post_Data = 8'h97; 
	12'h738 : Post_Data = 8'h97; 
	12'h739 : Post_Data = 8'h97; 
	12'h73A : Post_Data = 8'h97; 
	12'h73B : Post_Data = 8'h97; 
	12'h73C : Post_Data = 8'h97; 
	12'h73D : Post_Data = 8'h97; 
	12'h73E : Post_Data = 8'h97; 
	12'h73F : Post_Data = 8'h97; 
	12'h740 : Post_Data = 8'h97; 
	12'h741 : Post_Data = 8'h97; 
	12'h742 : Post_Data = 8'h97; 
	12'h743 : Post_Data = 8'h97; 
	12'h744 : Post_Data = 8'h97; 
	12'h745 : Post_Data = 8'h97; 
	12'h746 : Post_Data = 8'h97; 
	12'h747 : Post_Data = 8'h97; 
	12'h748 : Post_Data = 8'h98; 
	12'h749 : Post_Data = 8'h98; 
	12'h74A : Post_Data = 8'h98; 
	12'h74B : Post_Data = 8'h98; 
	12'h74C : Post_Data = 8'h98; 
	12'h74D : Post_Data = 8'h98; 
	12'h74E : Post_Data = 8'h98; 
	12'h74F : Post_Data = 8'h98; 
	12'h750 : Post_Data = 8'h98; 
	12'h751 : Post_Data = 8'h98; 
	12'h752 : Post_Data = 8'h98; 
	12'h753 : Post_Data = 8'h98; 
	12'h754 : Post_Data = 8'h98; 
	12'h755 : Post_Data = 8'h98; 
	12'h756 : Post_Data = 8'h98; 
	12'h757 : Post_Data = 8'h98; 
	12'h758 : Post_Data = 8'h98; 
	12'h759 : Post_Data = 8'h98; 
	12'h75A : Post_Data = 8'h98; 
	12'h75B : Post_Data = 8'h99; 
	12'h75C : Post_Data = 8'h99; 
	12'h75D : Post_Data = 8'h99; 
	12'h75E : Post_Data = 8'h99; 
	12'h75F : Post_Data = 8'h99; 
	12'h760 : Post_Data = 8'h99; 
	12'h761 : Post_Data = 8'h99; 
	12'h762 : Post_Data = 8'h99; 
	12'h763 : Post_Data = 8'h99; 
	12'h764 : Post_Data = 8'h99; 
	12'h765 : Post_Data = 8'h99; 
	12'h766 : Post_Data = 8'h99; 
	12'h767 : Post_Data = 8'h99; 
	12'h768 : Post_Data = 8'h99; 
	12'h769 : Post_Data = 8'h99; 
	12'h76A : Post_Data = 8'h99; 
	12'h76B : Post_Data = 8'h99; 
	12'h76C : Post_Data = 8'h99; 
	12'h76D : Post_Data = 8'h9A; 
	12'h76E : Post_Data = 8'h9A; 
	12'h76F : Post_Data = 8'h9A; 
	12'h770 : Post_Data = 8'h9A; 
	12'h771 : Post_Data = 8'h9A; 
	12'h772 : Post_Data = 8'h9A; 
	12'h773 : Post_Data = 8'h9A; 
	12'h774 : Post_Data = 8'h9A; 
	12'h775 : Post_Data = 8'h9A; 
	12'h776 : Post_Data = 8'h9A; 
	12'h777 : Post_Data = 8'h9A; 
	12'h778 : Post_Data = 8'h9A; 
	12'h779 : Post_Data = 8'h9A; 
	12'h77A : Post_Data = 8'h9A; 
	12'h77B : Post_Data = 8'h9A; 
	12'h77C : Post_Data = 8'h9A; 
	12'h77D : Post_Data = 8'h9A; 
	12'h77E : Post_Data = 8'h9A; 
	12'h77F : Post_Data = 8'h9A; 
	12'h780 : Post_Data = 8'h9B; 
	12'h781 : Post_Data = 8'h9B; 
	12'h782 : Post_Data = 8'h9B; 
	12'h783 : Post_Data = 8'h9B; 
	12'h784 : Post_Data = 8'h9B; 
	12'h785 : Post_Data = 8'h9B; 
	12'h786 : Post_Data = 8'h9B; 
	12'h787 : Post_Data = 8'h9B; 
	12'h788 : Post_Data = 8'h9B; 
	12'h789 : Post_Data = 8'h9B; 
	12'h78A : Post_Data = 8'h9B; 
	12'h78B : Post_Data = 8'h9B; 
	12'h78C : Post_Data = 8'h9B; 
	12'h78D : Post_Data = 8'h9B; 
	12'h78E : Post_Data = 8'h9B; 
	12'h78F : Post_Data = 8'h9B; 
	12'h790 : Post_Data = 8'h9B; 
	12'h791 : Post_Data = 8'h9B; 
	12'h792 : Post_Data = 8'h9B; 
	12'h793 : Post_Data = 8'h9C; 
	12'h794 : Post_Data = 8'h9C; 
	12'h795 : Post_Data = 8'h9C; 
	12'h796 : Post_Data = 8'h9C; 
	12'h797 : Post_Data = 8'h9C; 
	12'h798 : Post_Data = 8'h9C; 
	12'h799 : Post_Data = 8'h9C; 
	12'h79A : Post_Data = 8'h9C; 
	12'h79B : Post_Data = 8'h9C; 
	12'h79C : Post_Data = 8'h9C; 
	12'h79D : Post_Data = 8'h9C; 
	12'h79E : Post_Data = 8'h9C; 
	12'h79F : Post_Data = 8'h9C; 
	12'h7A0 : Post_Data = 8'h9C; 
	12'h7A1 : Post_Data = 8'h9C; 
	12'h7A2 : Post_Data = 8'h9C; 
	12'h7A3 : Post_Data = 8'h9C; 
	12'h7A4 : Post_Data = 8'h9C; 
	12'h7A5 : Post_Data = 8'h9D; 
	12'h7A6 : Post_Data = 8'h9D; 
	12'h7A7 : Post_Data = 8'h9D; 
	12'h7A8 : Post_Data = 8'h9D; 
	12'h7A9 : Post_Data = 8'h9D; 
	12'h7AA : Post_Data = 8'h9D; 
	12'h7AB : Post_Data = 8'h9D; 
	12'h7AC : Post_Data = 8'h9D; 
	12'h7AD : Post_Data = 8'h9D; 
	12'h7AE : Post_Data = 8'h9D; 
	12'h7AF : Post_Data = 8'h9D; 
	12'h7B0 : Post_Data = 8'h9D; 
	12'h7B1 : Post_Data = 8'h9D; 
	12'h7B2 : Post_Data = 8'h9D; 
	12'h7B3 : Post_Data = 8'h9D; 
	12'h7B4 : Post_Data = 8'h9D; 
	12'h7B5 : Post_Data = 8'h9D; 
	12'h7B6 : Post_Data = 8'h9D; 
	12'h7B7 : Post_Data = 8'h9D; 
	12'h7B8 : Post_Data = 8'h9E; 
	12'h7B9 : Post_Data = 8'h9E; 
	12'h7BA : Post_Data = 8'h9E; 
	12'h7BB : Post_Data = 8'h9E; 
	12'h7BC : Post_Data = 8'h9E; 
	12'h7BD : Post_Data = 8'h9E; 
	12'h7BE : Post_Data = 8'h9E; 
	12'h7BF : Post_Data = 8'h9E; 
	12'h7C0 : Post_Data = 8'h9E; 
	12'h7C1 : Post_Data = 8'h9E; 
	12'h7C2 : Post_Data = 8'h9E; 
	12'h7C3 : Post_Data = 8'h9E; 
	12'h7C4 : Post_Data = 8'h9E; 
	12'h7C5 : Post_Data = 8'h9E; 
	12'h7C6 : Post_Data = 8'h9E; 
	12'h7C7 : Post_Data = 8'h9E; 
	12'h7C8 : Post_Data = 8'h9E; 
	12'h7C9 : Post_Data = 8'h9E; 
	12'h7CA : Post_Data = 8'h9E; 
	12'h7CB : Post_Data = 8'h9F; 
	12'h7CC : Post_Data = 8'h9F; 
	12'h7CD : Post_Data = 8'h9F; 
	12'h7CE : Post_Data = 8'h9F; 
	12'h7CF : Post_Data = 8'h9F; 
	12'h7D0 : Post_Data = 8'h9F; 
	12'h7D1 : Post_Data = 8'h9F; 
	12'h7D2 : Post_Data = 8'h9F; 
	12'h7D3 : Post_Data = 8'h9F; 
	12'h7D4 : Post_Data = 8'h9F; 
	12'h7D5 : Post_Data = 8'h9F; 
	12'h7D6 : Post_Data = 8'h9F; 
	12'h7D7 : Post_Data = 8'h9F; 
	12'h7D8 : Post_Data = 8'h9F; 
	12'h7D9 : Post_Data = 8'h9F; 
	12'h7DA : Post_Data = 8'h9F; 
	12'h7DB : Post_Data = 8'h9F; 
	12'h7DC : Post_Data = 8'h9F; 
	12'h7DD : Post_Data = 8'h9F; 
	12'h7DE : Post_Data = 8'hA0; 
	12'h7DF : Post_Data = 8'hA0; 
	12'h7E0 : Post_Data = 8'hA0; 
	12'h7E1 : Post_Data = 8'hA0; 
	12'h7E2 : Post_Data = 8'hA0; 
	12'h7E3 : Post_Data = 8'hA0; 
	12'h7E4 : Post_Data = 8'hA0; 
	12'h7E5 : Post_Data = 8'hA0; 
	12'h7E6 : Post_Data = 8'hA0; 
	12'h7E7 : Post_Data = 8'hA0; 
	12'h7E8 : Post_Data = 8'hA0; 
	12'h7E9 : Post_Data = 8'hA0; 
	12'h7EA : Post_Data = 8'hA0; 
	12'h7EB : Post_Data = 8'hA0; 
	12'h7EC : Post_Data = 8'hA0; 
	12'h7ED : Post_Data = 8'hA0; 
	12'h7EE : Post_Data = 8'hA0; 
	12'h7EF : Post_Data = 8'hA0; 
	12'h7F0 : Post_Data = 8'hA0; 
	12'h7F1 : Post_Data = 8'hA1; 
	12'h7F2 : Post_Data = 8'hA1; 
	12'h7F3 : Post_Data = 8'hA1; 
	12'h7F4 : Post_Data = 8'hA1; 
	12'h7F5 : Post_Data = 8'hA1; 
	12'h7F6 : Post_Data = 8'hA1; 
	12'h7F7 : Post_Data = 8'hA1; 
	12'h7F8 : Post_Data = 8'hA1; 
	12'h7F9 : Post_Data = 8'hA1; 
	12'h7FA : Post_Data = 8'hA1; 
	12'h7FB : Post_Data = 8'hA1; 
	12'h7FC : Post_Data = 8'hA1; 
	12'h7FD : Post_Data = 8'hA1; 
	12'h7FE : Post_Data = 8'hA1; 
	12'h7FF : Post_Data = 8'hA1; 
	12'h800 : Post_Data = 8'hA1; 
	12'h801 : Post_Data = 8'hA1; 
	12'h802 : Post_Data = 8'hA1; 
	12'h803 : Post_Data = 8'hA1; 
	12'h804 : Post_Data = 8'hA2; 
	12'h805 : Post_Data = 8'hA2; 
	12'h806 : Post_Data = 8'hA2; 
	12'h807 : Post_Data = 8'hA2; 
	12'h808 : Post_Data = 8'hA2; 
	12'h809 : Post_Data = 8'hA2; 
	12'h80A : Post_Data = 8'hA2; 
	12'h80B : Post_Data = 8'hA2; 
	12'h80C : Post_Data = 8'hA2; 
	12'h80D : Post_Data = 8'hA2; 
	12'h80E : Post_Data = 8'hA2; 
	12'h80F : Post_Data = 8'hA2; 
	12'h810 : Post_Data = 8'hA2; 
	12'h811 : Post_Data = 8'hA2; 
	12'h812 : Post_Data = 8'hA2; 
	12'h813 : Post_Data = 8'hA2; 
	12'h814 : Post_Data = 8'hA2; 
	12'h815 : Post_Data = 8'hA2; 
	12'h816 : Post_Data = 8'hA2; 
	12'h817 : Post_Data = 8'hA3; 
	12'h818 : Post_Data = 8'hA3; 
	12'h819 : Post_Data = 8'hA3; 
	12'h81A : Post_Data = 8'hA3; 
	12'h81B : Post_Data = 8'hA3; 
	12'h81C : Post_Data = 8'hA3; 
	12'h81D : Post_Data = 8'hA3; 
	12'h81E : Post_Data = 8'hA3; 
	12'h81F : Post_Data = 8'hA3; 
	12'h820 : Post_Data = 8'hA3; 
	12'h821 : Post_Data = 8'hA3; 
	12'h822 : Post_Data = 8'hA3; 
	12'h823 : Post_Data = 8'hA3; 
	12'h824 : Post_Data = 8'hA3; 
	12'h825 : Post_Data = 8'hA3; 
	12'h826 : Post_Data = 8'hA3; 
	12'h827 : Post_Data = 8'hA3; 
	12'h828 : Post_Data = 8'hA3; 
	12'h829 : Post_Data = 8'hA3; 
	12'h82A : Post_Data = 8'hA4; 
	12'h82B : Post_Data = 8'hA4; 
	12'h82C : Post_Data = 8'hA4; 
	12'h82D : Post_Data = 8'hA4; 
	12'h82E : Post_Data = 8'hA4; 
	12'h82F : Post_Data = 8'hA4; 
	12'h830 : Post_Data = 8'hA4; 
	12'h831 : Post_Data = 8'hA4; 
	12'h832 : Post_Data = 8'hA4; 
	12'h833 : Post_Data = 8'hA4; 
	12'h834 : Post_Data = 8'hA4; 
	12'h835 : Post_Data = 8'hA4; 
	12'h836 : Post_Data = 8'hA4; 
	12'h837 : Post_Data = 8'hA4; 
	12'h838 : Post_Data = 8'hA4; 
	12'h839 : Post_Data = 8'hA4; 
	12'h83A : Post_Data = 8'hA4; 
	12'h83B : Post_Data = 8'hA4; 
	12'h83C : Post_Data = 8'hA4; 
	12'h83D : Post_Data = 8'hA5; 
	12'h83E : Post_Data = 8'hA5; 
	12'h83F : Post_Data = 8'hA5; 
	12'h840 : Post_Data = 8'hA5; 
	12'h841 : Post_Data = 8'hA5; 
	12'h842 : Post_Data = 8'hA5; 
	12'h843 : Post_Data = 8'hA5; 
	12'h844 : Post_Data = 8'hA5; 
	12'h845 : Post_Data = 8'hA5; 
	12'h846 : Post_Data = 8'hA5; 
	12'h847 : Post_Data = 8'hA5; 
	12'h848 : Post_Data = 8'hA5; 
	12'h849 : Post_Data = 8'hA5; 
	12'h84A : Post_Data = 8'hA5; 
	12'h84B : Post_Data = 8'hA5; 
	12'h84C : Post_Data = 8'hA5; 
	12'h84D : Post_Data = 8'hA5; 
	12'h84E : Post_Data = 8'hA5; 
	12'h84F : Post_Data = 8'hA5; 
	12'h850 : Post_Data = 8'hA5; 
	12'h851 : Post_Data = 8'hA6; 
	12'h852 : Post_Data = 8'hA6; 
	12'h853 : Post_Data = 8'hA6; 
	12'h854 : Post_Data = 8'hA6; 
	12'h855 : Post_Data = 8'hA6; 
	12'h856 : Post_Data = 8'hA6; 
	12'h857 : Post_Data = 8'hA6; 
	12'h858 : Post_Data = 8'hA6; 
	12'h859 : Post_Data = 8'hA6; 
	12'h85A : Post_Data = 8'hA6; 
	12'h85B : Post_Data = 8'hA6; 
	12'h85C : Post_Data = 8'hA6; 
	12'h85D : Post_Data = 8'hA6; 
	12'h85E : Post_Data = 8'hA6; 
	12'h85F : Post_Data = 8'hA6; 
	12'h860 : Post_Data = 8'hA6; 
	12'h861 : Post_Data = 8'hA6; 
	12'h862 : Post_Data = 8'hA6; 
	12'h863 : Post_Data = 8'hA6; 
	12'h864 : Post_Data = 8'hA7; 
	12'h865 : Post_Data = 8'hA7; 
	12'h866 : Post_Data = 8'hA7; 
	12'h867 : Post_Data = 8'hA7; 
	12'h868 : Post_Data = 8'hA7; 
	12'h869 : Post_Data = 8'hA7; 
	12'h86A : Post_Data = 8'hA7; 
	12'h86B : Post_Data = 8'hA7; 
	12'h86C : Post_Data = 8'hA7; 
	12'h86D : Post_Data = 8'hA7; 
	12'h86E : Post_Data = 8'hA7; 
	12'h86F : Post_Data = 8'hA7; 
	12'h870 : Post_Data = 8'hA7; 
	12'h871 : Post_Data = 8'hA7; 
	12'h872 : Post_Data = 8'hA7; 
	12'h873 : Post_Data = 8'hA7; 
	12'h874 : Post_Data = 8'hA7; 
	12'h875 : Post_Data = 8'hA7; 
	12'h876 : Post_Data = 8'hA7; 
	12'h877 : Post_Data = 8'hA8; 
	12'h878 : Post_Data = 8'hA8; 
	12'h879 : Post_Data = 8'hA8; 
	12'h87A : Post_Data = 8'hA8; 
	12'h87B : Post_Data = 8'hA8; 
	12'h87C : Post_Data = 8'hA8; 
	12'h87D : Post_Data = 8'hA8; 
	12'h87E : Post_Data = 8'hA8; 
	12'h87F : Post_Data = 8'hA8; 
	12'h880 : Post_Data = 8'hA8; 
	12'h881 : Post_Data = 8'hA8; 
	12'h882 : Post_Data = 8'hA8; 
	12'h883 : Post_Data = 8'hA8; 
	12'h884 : Post_Data = 8'hA8; 
	12'h885 : Post_Data = 8'hA8; 
	12'h886 : Post_Data = 8'hA8; 
	12'h887 : Post_Data = 8'hA8; 
	12'h888 : Post_Data = 8'hA8; 
	12'h889 : Post_Data = 8'hA8; 
	12'h88A : Post_Data = 8'hA8; 
	12'h88B : Post_Data = 8'hA9; 
	12'h88C : Post_Data = 8'hA9; 
	12'h88D : Post_Data = 8'hA9; 
	12'h88E : Post_Data = 8'hA9; 
	12'h88F : Post_Data = 8'hA9; 
	12'h890 : Post_Data = 8'hA9; 
	12'h891 : Post_Data = 8'hA9; 
	12'h892 : Post_Data = 8'hA9; 
	12'h893 : Post_Data = 8'hA9; 
	12'h894 : Post_Data = 8'hA9; 
	12'h895 : Post_Data = 8'hA9; 
	12'h896 : Post_Data = 8'hA9; 
	12'h897 : Post_Data = 8'hA9; 
	12'h898 : Post_Data = 8'hA9; 
	12'h899 : Post_Data = 8'hA9; 
	12'h89A : Post_Data = 8'hA9; 
	12'h89B : Post_Data = 8'hA9; 
	12'h89C : Post_Data = 8'hA9; 
	12'h89D : Post_Data = 8'hA9; 
	12'h89E : Post_Data = 8'hAA; 
	12'h89F : Post_Data = 8'hAA; 
	12'h8A0 : Post_Data = 8'hAA; 
	12'h8A1 : Post_Data = 8'hAA; 
	12'h8A2 : Post_Data = 8'hAA; 
	12'h8A3 : Post_Data = 8'hAA; 
	12'h8A4 : Post_Data = 8'hAA; 
	12'h8A5 : Post_Data = 8'hAA; 
	12'h8A6 : Post_Data = 8'hAA; 
	12'h8A7 : Post_Data = 8'hAA; 
	12'h8A8 : Post_Data = 8'hAA; 
	12'h8A9 : Post_Data = 8'hAA; 
	12'h8AA : Post_Data = 8'hAA; 
	12'h8AB : Post_Data = 8'hAA; 
	12'h8AC : Post_Data = 8'hAA; 
	12'h8AD : Post_Data = 8'hAA; 
	12'h8AE : Post_Data = 8'hAA; 
	12'h8AF : Post_Data = 8'hAA; 
	12'h8B0 : Post_Data = 8'hAA; 
	12'h8B1 : Post_Data = 8'hAA; 
	12'h8B2 : Post_Data = 8'hAB; 
	12'h8B3 : Post_Data = 8'hAB; 
	12'h8B4 : Post_Data = 8'hAB; 
	12'h8B5 : Post_Data = 8'hAB; 
	12'h8B6 : Post_Data = 8'hAB; 
	12'h8B7 : Post_Data = 8'hAB; 
	12'h8B8 : Post_Data = 8'hAB; 
	12'h8B9 : Post_Data = 8'hAB; 
	12'h8BA : Post_Data = 8'hAB; 
	12'h8BB : Post_Data = 8'hAB; 
	12'h8BC : Post_Data = 8'hAB; 
	12'h8BD : Post_Data = 8'hAB; 
	12'h8BE : Post_Data = 8'hAB; 
	12'h8BF : Post_Data = 8'hAB; 
	12'h8C0 : Post_Data = 8'hAB; 
	12'h8C1 : Post_Data = 8'hAB; 
	12'h8C2 : Post_Data = 8'hAB; 
	12'h8C3 : Post_Data = 8'hAB; 
	12'h8C4 : Post_Data = 8'hAB; 
	12'h8C5 : Post_Data = 8'hAC; 
	12'h8C6 : Post_Data = 8'hAC; 
	12'h8C7 : Post_Data = 8'hAC; 
	12'h8C8 : Post_Data = 8'hAC; 
	12'h8C9 : Post_Data = 8'hAC; 
	12'h8CA : Post_Data = 8'hAC; 
	12'h8CB : Post_Data = 8'hAC; 
	12'h8CC : Post_Data = 8'hAC; 
	12'h8CD : Post_Data = 8'hAC; 
	12'h8CE : Post_Data = 8'hAC; 
	12'h8CF : Post_Data = 8'hAC; 
	12'h8D0 : Post_Data = 8'hAC; 
	12'h8D1 : Post_Data = 8'hAC; 
	12'h8D2 : Post_Data = 8'hAC; 
	12'h8D3 : Post_Data = 8'hAC; 
	12'h8D4 : Post_Data = 8'hAC; 
	12'h8D5 : Post_Data = 8'hAC; 
	12'h8D6 : Post_Data = 8'hAC; 
	12'h8D7 : Post_Data = 8'hAC; 
	12'h8D8 : Post_Data = 8'hAC; 
	12'h8D9 : Post_Data = 8'hAD; 
	12'h8DA : Post_Data = 8'hAD; 
	12'h8DB : Post_Data = 8'hAD; 
	12'h8DC : Post_Data = 8'hAD; 
	12'h8DD : Post_Data = 8'hAD; 
	12'h8DE : Post_Data = 8'hAD; 
	12'h8DF : Post_Data = 8'hAD; 
	12'h8E0 : Post_Data = 8'hAD; 
	12'h8E1 : Post_Data = 8'hAD; 
	12'h8E2 : Post_Data = 8'hAD; 
	12'h8E3 : Post_Data = 8'hAD; 
	12'h8E4 : Post_Data = 8'hAD; 
	12'h8E5 : Post_Data = 8'hAD; 
	12'h8E6 : Post_Data = 8'hAD; 
	12'h8E7 : Post_Data = 8'hAD; 
	12'h8E8 : Post_Data = 8'hAD; 
	12'h8E9 : Post_Data = 8'hAD; 
	12'h8EA : Post_Data = 8'hAD; 
	12'h8EB : Post_Data = 8'hAD; 
	12'h8EC : Post_Data = 8'hAD; 
	12'h8ED : Post_Data = 8'hAE; 
	12'h8EE : Post_Data = 8'hAE; 
	12'h8EF : Post_Data = 8'hAE; 
	12'h8F0 : Post_Data = 8'hAE; 
	12'h8F1 : Post_Data = 8'hAE; 
	12'h8F2 : Post_Data = 8'hAE; 
	12'h8F3 : Post_Data = 8'hAE; 
	12'h8F4 : Post_Data = 8'hAE; 
	12'h8F5 : Post_Data = 8'hAE; 
	12'h8F6 : Post_Data = 8'hAE; 
	12'h8F7 : Post_Data = 8'hAE; 
	12'h8F8 : Post_Data = 8'hAE; 
	12'h8F9 : Post_Data = 8'hAE; 
	12'h8FA : Post_Data = 8'hAE; 
	12'h8FB : Post_Data = 8'hAE; 
	12'h8FC : Post_Data = 8'hAE; 
	12'h8FD : Post_Data = 8'hAE; 
	12'h8FE : Post_Data = 8'hAE; 
	12'h8FF : Post_Data = 8'hAE; 
	12'h900 : Post_Data = 8'hAE; 
	12'h901 : Post_Data = 8'hAF; 
	12'h902 : Post_Data = 8'hAF; 
	12'h903 : Post_Data = 8'hAF; 
	12'h904 : Post_Data = 8'hAF; 
	12'h905 : Post_Data = 8'hAF; 
	12'h906 : Post_Data = 8'hAF; 
	12'h907 : Post_Data = 8'hAF; 
	12'h908 : Post_Data = 8'hAF; 
	12'h909 : Post_Data = 8'hAF; 
	12'h90A : Post_Data = 8'hAF; 
	12'h90B : Post_Data = 8'hAF; 
	12'h90C : Post_Data = 8'hAF; 
	12'h90D : Post_Data = 8'hAF; 
	12'h90E : Post_Data = 8'hAF; 
	12'h90F : Post_Data = 8'hAF; 
	12'h910 : Post_Data = 8'hAF; 
	12'h911 : Post_Data = 8'hAF; 
	12'h912 : Post_Data = 8'hAF; 
	12'h913 : Post_Data = 8'hAF; 
	12'h914 : Post_Data = 8'hB0; 
	12'h915 : Post_Data = 8'hB0; 
	12'h916 : Post_Data = 8'hB0; 
	12'h917 : Post_Data = 8'hB0; 
	12'h918 : Post_Data = 8'hB0; 
	12'h919 : Post_Data = 8'hB0; 
	12'h91A : Post_Data = 8'hB0; 
	12'h91B : Post_Data = 8'hB0; 
	12'h91C : Post_Data = 8'hB0; 
	12'h91D : Post_Data = 8'hB0; 
	12'h91E : Post_Data = 8'hB0; 
	12'h91F : Post_Data = 8'hB0; 
	12'h920 : Post_Data = 8'hB0; 
	12'h921 : Post_Data = 8'hB0; 
	12'h922 : Post_Data = 8'hB0; 
	12'h923 : Post_Data = 8'hB0; 
	12'h924 : Post_Data = 8'hB0; 
	12'h925 : Post_Data = 8'hB0; 
	12'h926 : Post_Data = 8'hB0; 
	12'h927 : Post_Data = 8'hB0; 
	12'h928 : Post_Data = 8'hB1; 
	12'h929 : Post_Data = 8'hB1; 
	12'h92A : Post_Data = 8'hB1; 
	12'h92B : Post_Data = 8'hB1; 
	12'h92C : Post_Data = 8'hB1; 
	12'h92D : Post_Data = 8'hB1; 
	12'h92E : Post_Data = 8'hB1; 
	12'h92F : Post_Data = 8'hB1; 
	12'h930 : Post_Data = 8'hB1; 
	12'h931 : Post_Data = 8'hB1; 
	12'h932 : Post_Data = 8'hB1; 
	12'h933 : Post_Data = 8'hB1; 
	12'h934 : Post_Data = 8'hB1; 
	12'h935 : Post_Data = 8'hB1; 
	12'h936 : Post_Data = 8'hB1; 
	12'h937 : Post_Data = 8'hB1; 
	12'h938 : Post_Data = 8'hB1; 
	12'h939 : Post_Data = 8'hB1; 
	12'h93A : Post_Data = 8'hB1; 
	12'h93B : Post_Data = 8'hB1; 
	12'h93C : Post_Data = 8'hB2; 
	12'h93D : Post_Data = 8'hB2; 
	12'h93E : Post_Data = 8'hB2; 
	12'h93F : Post_Data = 8'hB2; 
	12'h940 : Post_Data = 8'hB2; 
	12'h941 : Post_Data = 8'hB2; 
	12'h942 : Post_Data = 8'hB2; 
	12'h943 : Post_Data = 8'hB2; 
	12'h944 : Post_Data = 8'hB2; 
	12'h945 : Post_Data = 8'hB2; 
	12'h946 : Post_Data = 8'hB2; 
	12'h947 : Post_Data = 8'hB2; 
	12'h948 : Post_Data = 8'hB2; 
	12'h949 : Post_Data = 8'hB2; 
	12'h94A : Post_Data = 8'hB2; 
	12'h94B : Post_Data = 8'hB2; 
	12'h94C : Post_Data = 8'hB2; 
	12'h94D : Post_Data = 8'hB2; 
	12'h94E : Post_Data = 8'hB2; 
	12'h94F : Post_Data = 8'hB2; 
	12'h950 : Post_Data = 8'hB3; 
	12'h951 : Post_Data = 8'hB3; 
	12'h952 : Post_Data = 8'hB3; 
	12'h953 : Post_Data = 8'hB3; 
	12'h954 : Post_Data = 8'hB3; 
	12'h955 : Post_Data = 8'hB3; 
	12'h956 : Post_Data = 8'hB3; 
	12'h957 : Post_Data = 8'hB3; 
	12'h958 : Post_Data = 8'hB3; 
	12'h959 : Post_Data = 8'hB3; 
	12'h95A : Post_Data = 8'hB3; 
	12'h95B : Post_Data = 8'hB3; 
	12'h95C : Post_Data = 8'hB3; 
	12'h95D : Post_Data = 8'hB3; 
	12'h95E : Post_Data = 8'hB3; 
	12'h95F : Post_Data = 8'hB3; 
	12'h960 : Post_Data = 8'hB3; 
	12'h961 : Post_Data = 8'hB3; 
	12'h962 : Post_Data = 8'hB3; 
	12'h963 : Post_Data = 8'hB3; 
	12'h964 : Post_Data = 8'hB4; 
	12'h965 : Post_Data = 8'hB4; 
	12'h966 : Post_Data = 8'hB4; 
	12'h967 : Post_Data = 8'hB4; 
	12'h968 : Post_Data = 8'hB4; 
	12'h969 : Post_Data = 8'hB4; 
	12'h96A : Post_Data = 8'hB4; 
	12'h96B : Post_Data = 8'hB4; 
	12'h96C : Post_Data = 8'hB4; 
	12'h96D : Post_Data = 8'hB4; 
	12'h96E : Post_Data = 8'hB4; 
	12'h96F : Post_Data = 8'hB4; 
	12'h970 : Post_Data = 8'hB4; 
	12'h971 : Post_Data = 8'hB4; 
	12'h972 : Post_Data = 8'hB4; 
	12'h973 : Post_Data = 8'hB4; 
	12'h974 : Post_Data = 8'hB4; 
	12'h975 : Post_Data = 8'hB4; 
	12'h976 : Post_Data = 8'hB4; 
	12'h977 : Post_Data = 8'hB4; 
	12'h978 : Post_Data = 8'hB4; 
	12'h979 : Post_Data = 8'hB5; 
	12'h97A : Post_Data = 8'hB5; 
	12'h97B : Post_Data = 8'hB5; 
	12'h97C : Post_Data = 8'hB5; 
	12'h97D : Post_Data = 8'hB5; 
	12'h97E : Post_Data = 8'hB5; 
	12'h97F : Post_Data = 8'hB5; 
	12'h980 : Post_Data = 8'hB5; 
	12'h981 : Post_Data = 8'hB5; 
	12'h982 : Post_Data = 8'hB5; 
	12'h983 : Post_Data = 8'hB5; 
	12'h984 : Post_Data = 8'hB5; 
	12'h985 : Post_Data = 8'hB5; 
	12'h986 : Post_Data = 8'hB5; 
	12'h987 : Post_Data = 8'hB5; 
	12'h988 : Post_Data = 8'hB5; 
	12'h989 : Post_Data = 8'hB5; 
	12'h98A : Post_Data = 8'hB5; 
	12'h98B : Post_Data = 8'hB5; 
	12'h98C : Post_Data = 8'hB5; 
	12'h98D : Post_Data = 8'hB6; 
	12'h98E : Post_Data = 8'hB6; 
	12'h98F : Post_Data = 8'hB6; 
	12'h990 : Post_Data = 8'hB6; 
	12'h991 : Post_Data = 8'hB6; 
	12'h992 : Post_Data = 8'hB6; 
	12'h993 : Post_Data = 8'hB6; 
	12'h994 : Post_Data = 8'hB6; 
	12'h995 : Post_Data = 8'hB6; 
	12'h996 : Post_Data = 8'hB6; 
	12'h997 : Post_Data = 8'hB6; 
	12'h998 : Post_Data = 8'hB6; 
	12'h999 : Post_Data = 8'hB6; 
	12'h99A : Post_Data = 8'hB6; 
	12'h99B : Post_Data = 8'hB6; 
	12'h99C : Post_Data = 8'hB6; 
	12'h99D : Post_Data = 8'hB6; 
	12'h99E : Post_Data = 8'hB6; 
	12'h99F : Post_Data = 8'hB6; 
	12'h9A0 : Post_Data = 8'hB6; 
	12'h9A1 : Post_Data = 8'hB7; 
	12'h9A2 : Post_Data = 8'hB7; 
	12'h9A3 : Post_Data = 8'hB7; 
	12'h9A4 : Post_Data = 8'hB7; 
	12'h9A5 : Post_Data = 8'hB7; 
	12'h9A6 : Post_Data = 8'hB7; 
	12'h9A7 : Post_Data = 8'hB7; 
	12'h9A8 : Post_Data = 8'hB7; 
	12'h9A9 : Post_Data = 8'hB7; 
	12'h9AA : Post_Data = 8'hB7; 
	12'h9AB : Post_Data = 8'hB7; 
	12'h9AC : Post_Data = 8'hB7; 
	12'h9AD : Post_Data = 8'hB7; 
	12'h9AE : Post_Data = 8'hB7; 
	12'h9AF : Post_Data = 8'hB7; 
	12'h9B0 : Post_Data = 8'hB7; 
	12'h9B1 : Post_Data = 8'hB7; 
	12'h9B2 : Post_Data = 8'hB7; 
	12'h9B3 : Post_Data = 8'hB7; 
	12'h9B4 : Post_Data = 8'hB7; 
	12'h9B5 : Post_Data = 8'hB8; 
	12'h9B6 : Post_Data = 8'hB8; 
	12'h9B7 : Post_Data = 8'hB8; 
	12'h9B8 : Post_Data = 8'hB8; 
	12'h9B9 : Post_Data = 8'hB8; 
	12'h9BA : Post_Data = 8'hB8; 
	12'h9BB : Post_Data = 8'hB8; 
	12'h9BC : Post_Data = 8'hB8; 
	12'h9BD : Post_Data = 8'hB8; 
	12'h9BE : Post_Data = 8'hB8; 
	12'h9BF : Post_Data = 8'hB8; 
	12'h9C0 : Post_Data = 8'hB8; 
	12'h9C1 : Post_Data = 8'hB8; 
	12'h9C2 : Post_Data = 8'hB8; 
	12'h9C3 : Post_Data = 8'hB8; 
	12'h9C4 : Post_Data = 8'hB8; 
	12'h9C5 : Post_Data = 8'hB8; 
	12'h9C6 : Post_Data = 8'hB8; 
	12'h9C7 : Post_Data = 8'hB8; 
	12'h9C8 : Post_Data = 8'hB8; 
	12'h9C9 : Post_Data = 8'hB8; 
	12'h9CA : Post_Data = 8'hB9; 
	12'h9CB : Post_Data = 8'hB9; 
	12'h9CC : Post_Data = 8'hB9; 
	12'h9CD : Post_Data = 8'hB9; 
	12'h9CE : Post_Data = 8'hB9; 
	12'h9CF : Post_Data = 8'hB9; 
	12'h9D0 : Post_Data = 8'hB9; 
	12'h9D1 : Post_Data = 8'hB9; 
	12'h9D2 : Post_Data = 8'hB9; 
	12'h9D3 : Post_Data = 8'hB9; 
	12'h9D4 : Post_Data = 8'hB9; 
	12'h9D5 : Post_Data = 8'hB9; 
	12'h9D6 : Post_Data = 8'hB9; 
	12'h9D7 : Post_Data = 8'hB9; 
	12'h9D8 : Post_Data = 8'hB9; 
	12'h9D9 : Post_Data = 8'hB9; 
	12'h9DA : Post_Data = 8'hB9; 
	12'h9DB : Post_Data = 8'hB9; 
	12'h9DC : Post_Data = 8'hB9; 
	12'h9DD : Post_Data = 8'hB9; 
	12'h9DE : Post_Data = 8'hBA; 
	12'h9DF : Post_Data = 8'hBA; 
	12'h9E0 : Post_Data = 8'hBA; 
	12'h9E1 : Post_Data = 8'hBA; 
	12'h9E2 : Post_Data = 8'hBA; 
	12'h9E3 : Post_Data = 8'hBA; 
	12'h9E4 : Post_Data = 8'hBA; 
	12'h9E5 : Post_Data = 8'hBA; 
	12'h9E6 : Post_Data = 8'hBA; 
	12'h9E7 : Post_Data = 8'hBA; 
	12'h9E8 : Post_Data = 8'hBA; 
	12'h9E9 : Post_Data = 8'hBA; 
	12'h9EA : Post_Data = 8'hBA; 
	12'h9EB : Post_Data = 8'hBA; 
	12'h9EC : Post_Data = 8'hBA; 
	12'h9ED : Post_Data = 8'hBA; 
	12'h9EE : Post_Data = 8'hBA; 
	12'h9EF : Post_Data = 8'hBA; 
	12'h9F0 : Post_Data = 8'hBA; 
	12'h9F1 : Post_Data = 8'hBA; 
	12'h9F2 : Post_Data = 8'hBB; 
	12'h9F3 : Post_Data = 8'hBB; 
	12'h9F4 : Post_Data = 8'hBB; 
	12'h9F5 : Post_Data = 8'hBB; 
	12'h9F6 : Post_Data = 8'hBB; 
	12'h9F7 : Post_Data = 8'hBB; 
	12'h9F8 : Post_Data = 8'hBB; 
	12'h9F9 : Post_Data = 8'hBB; 
	12'h9FA : Post_Data = 8'hBB; 
	12'h9FB : Post_Data = 8'hBB; 
	12'h9FC : Post_Data = 8'hBB; 
	12'h9FD : Post_Data = 8'hBB; 
	12'h9FE : Post_Data = 8'hBB; 
	12'h9FF : Post_Data = 8'hBB; 
	12'hA00 : Post_Data = 8'hBB; 
	12'hA01 : Post_Data = 8'hBB; 
	12'hA02 : Post_Data = 8'hBB; 
	12'hA03 : Post_Data = 8'hBB; 
	12'hA04 : Post_Data = 8'hBB; 
	12'hA05 : Post_Data = 8'hBB; 
	12'hA06 : Post_Data = 8'hBB; 
	12'hA07 : Post_Data = 8'hBC; 
	12'hA08 : Post_Data = 8'hBC; 
	12'hA09 : Post_Data = 8'hBC; 
	12'hA0A : Post_Data = 8'hBC; 
	12'hA0B : Post_Data = 8'hBC; 
	12'hA0C : Post_Data = 8'hBC; 
	12'hA0D : Post_Data = 8'hBC; 
	12'hA0E : Post_Data = 8'hBC; 
	12'hA0F : Post_Data = 8'hBC; 
	12'hA10 : Post_Data = 8'hBC; 
	12'hA11 : Post_Data = 8'hBC; 
	12'hA12 : Post_Data = 8'hBC; 
	12'hA13 : Post_Data = 8'hBC; 
	12'hA14 : Post_Data = 8'hBC; 
	12'hA15 : Post_Data = 8'hBC; 
	12'hA16 : Post_Data = 8'hBC; 
	12'hA17 : Post_Data = 8'hBC; 
	12'hA18 : Post_Data = 8'hBC; 
	12'hA19 : Post_Data = 8'hBC; 
	12'hA1A : Post_Data = 8'hBC; 
	12'hA1B : Post_Data = 8'hBC; 
	12'hA1C : Post_Data = 8'hBD; 
	12'hA1D : Post_Data = 8'hBD; 
	12'hA1E : Post_Data = 8'hBD; 
	12'hA1F : Post_Data = 8'hBD; 
	12'hA20 : Post_Data = 8'hBD; 
	12'hA21 : Post_Data = 8'hBD; 
	12'hA22 : Post_Data = 8'hBD; 
	12'hA23 : Post_Data = 8'hBD; 
	12'hA24 : Post_Data = 8'hBD; 
	12'hA25 : Post_Data = 8'hBD; 
	12'hA26 : Post_Data = 8'hBD; 
	12'hA27 : Post_Data = 8'hBD; 
	12'hA28 : Post_Data = 8'hBD; 
	12'hA29 : Post_Data = 8'hBD; 
	12'hA2A : Post_Data = 8'hBD; 
	12'hA2B : Post_Data = 8'hBD; 
	12'hA2C : Post_Data = 8'hBD; 
	12'hA2D : Post_Data = 8'hBD; 
	12'hA2E : Post_Data = 8'hBD; 
	12'hA2F : Post_Data = 8'hBD; 
	12'hA30 : Post_Data = 8'hBE; 
	12'hA31 : Post_Data = 8'hBE; 
	12'hA32 : Post_Data = 8'hBE; 
	12'hA33 : Post_Data = 8'hBE; 
	12'hA34 : Post_Data = 8'hBE; 
	12'hA35 : Post_Data = 8'hBE; 
	12'hA36 : Post_Data = 8'hBE; 
	12'hA37 : Post_Data = 8'hBE; 
	12'hA38 : Post_Data = 8'hBE; 
	12'hA39 : Post_Data = 8'hBE; 
	12'hA3A : Post_Data = 8'hBE; 
	12'hA3B : Post_Data = 8'hBE; 
	12'hA3C : Post_Data = 8'hBE; 
	12'hA3D : Post_Data = 8'hBE; 
	12'hA3E : Post_Data = 8'hBE; 
	12'hA3F : Post_Data = 8'hBE; 
	12'hA40 : Post_Data = 8'hBE; 
	12'hA41 : Post_Data = 8'hBE; 
	12'hA42 : Post_Data = 8'hBE; 
	12'hA43 : Post_Data = 8'hBE; 
	12'hA44 : Post_Data = 8'hBE; 
	12'hA45 : Post_Data = 8'hBF; 
	12'hA46 : Post_Data = 8'hBF; 
	12'hA47 : Post_Data = 8'hBF; 
	12'hA48 : Post_Data = 8'hBF; 
	12'hA49 : Post_Data = 8'hBF; 
	12'hA4A : Post_Data = 8'hBF; 
	12'hA4B : Post_Data = 8'hBF; 
	12'hA4C : Post_Data = 8'hBF; 
	12'hA4D : Post_Data = 8'hBF; 
	12'hA4E : Post_Data = 8'hBF; 
	12'hA4F : Post_Data = 8'hBF; 
	12'hA50 : Post_Data = 8'hBF; 
	12'hA51 : Post_Data = 8'hBF; 
	12'hA52 : Post_Data = 8'hBF; 
	12'hA53 : Post_Data = 8'hBF; 
	12'hA54 : Post_Data = 8'hBF; 
	12'hA55 : Post_Data = 8'hBF; 
	12'hA56 : Post_Data = 8'hBF; 
	12'hA57 : Post_Data = 8'hBF; 
	12'hA58 : Post_Data = 8'hBF; 
	12'hA59 : Post_Data = 8'hBF; 
	12'hA5A : Post_Data = 8'hC0; 
	12'hA5B : Post_Data = 8'hC0; 
	12'hA5C : Post_Data = 8'hC0; 
	12'hA5D : Post_Data = 8'hC0; 
	12'hA5E : Post_Data = 8'hC0; 
	12'hA5F : Post_Data = 8'hC0; 
	12'hA60 : Post_Data = 8'hC0; 
	12'hA61 : Post_Data = 8'hC0; 
	12'hA62 : Post_Data = 8'hC0; 
	12'hA63 : Post_Data = 8'hC0; 
	12'hA64 : Post_Data = 8'hC0; 
	12'hA65 : Post_Data = 8'hC0; 
	12'hA66 : Post_Data = 8'hC0; 
	12'hA67 : Post_Data = 8'hC0; 
	12'hA68 : Post_Data = 8'hC0; 
	12'hA69 : Post_Data = 8'hC0; 
	12'hA6A : Post_Data = 8'hC0; 
	12'hA6B : Post_Data = 8'hC0; 
	12'hA6C : Post_Data = 8'hC0; 
	12'hA6D : Post_Data = 8'hC0; 
	12'hA6E : Post_Data = 8'hC1; 
	12'hA6F : Post_Data = 8'hC1; 
	12'hA70 : Post_Data = 8'hC1; 
	12'hA71 : Post_Data = 8'hC1; 
	12'hA72 : Post_Data = 8'hC1; 
	12'hA73 : Post_Data = 8'hC1; 
	12'hA74 : Post_Data = 8'hC1; 
	12'hA75 : Post_Data = 8'hC1; 
	12'hA76 : Post_Data = 8'hC1; 
	12'hA77 : Post_Data = 8'hC1; 
	12'hA78 : Post_Data = 8'hC1; 
	12'hA79 : Post_Data = 8'hC1; 
	12'hA7A : Post_Data = 8'hC1; 
	12'hA7B : Post_Data = 8'hC1; 
	12'hA7C : Post_Data = 8'hC1; 
	12'hA7D : Post_Data = 8'hC1; 
	12'hA7E : Post_Data = 8'hC1; 
	12'hA7F : Post_Data = 8'hC1; 
	12'hA80 : Post_Data = 8'hC1; 
	12'hA81 : Post_Data = 8'hC1; 
	12'hA82 : Post_Data = 8'hC1; 
	12'hA83 : Post_Data = 8'hC2; 
	12'hA84 : Post_Data = 8'hC2; 
	12'hA85 : Post_Data = 8'hC2; 
	12'hA86 : Post_Data = 8'hC2; 
	12'hA87 : Post_Data = 8'hC2; 
	12'hA88 : Post_Data = 8'hC2; 
	12'hA89 : Post_Data = 8'hC2; 
	12'hA8A : Post_Data = 8'hC2; 
	12'hA8B : Post_Data = 8'hC2; 
	12'hA8C : Post_Data = 8'hC2; 
	12'hA8D : Post_Data = 8'hC2; 
	12'hA8E : Post_Data = 8'hC2; 
	12'hA8F : Post_Data = 8'hC2; 
	12'hA90 : Post_Data = 8'hC2; 
	12'hA91 : Post_Data = 8'hC2; 
	12'hA92 : Post_Data = 8'hC2; 
	12'hA93 : Post_Data = 8'hC2; 
	12'hA94 : Post_Data = 8'hC2; 
	12'hA95 : Post_Data = 8'hC2; 
	12'hA96 : Post_Data = 8'hC2; 
	12'hA97 : Post_Data = 8'hC2; 
	12'hA98 : Post_Data = 8'hC3; 
	12'hA99 : Post_Data = 8'hC3; 
	12'hA9A : Post_Data = 8'hC3; 
	12'hA9B : Post_Data = 8'hC3; 
	12'hA9C : Post_Data = 8'hC3; 
	12'hA9D : Post_Data = 8'hC3; 
	12'hA9E : Post_Data = 8'hC3; 
	12'hA9F : Post_Data = 8'hC3; 
	12'hAA0 : Post_Data = 8'hC3; 
	12'hAA1 : Post_Data = 8'hC3; 
	12'hAA2 : Post_Data = 8'hC3; 
	12'hAA3 : Post_Data = 8'hC3; 
	12'hAA4 : Post_Data = 8'hC3; 
	12'hAA5 : Post_Data = 8'hC3; 
	12'hAA6 : Post_Data = 8'hC3; 
	12'hAA7 : Post_Data = 8'hC3; 
	12'hAA8 : Post_Data = 8'hC3; 
	12'hAA9 : Post_Data = 8'hC3; 
	12'hAAA : Post_Data = 8'hC3; 
	12'hAAB : Post_Data = 8'hC3; 
	12'hAAC : Post_Data = 8'hC3; 
	12'hAAD : Post_Data = 8'hC4; 
	12'hAAE : Post_Data = 8'hC4; 
	12'hAAF : Post_Data = 8'hC4; 
	12'hAB0 : Post_Data = 8'hC4; 
	12'hAB1 : Post_Data = 8'hC4; 
	12'hAB2 : Post_Data = 8'hC4; 
	12'hAB3 : Post_Data = 8'hC4; 
	12'hAB4 : Post_Data = 8'hC4; 
	12'hAB5 : Post_Data = 8'hC4; 
	12'hAB6 : Post_Data = 8'hC4; 
	12'hAB7 : Post_Data = 8'hC4; 
	12'hAB8 : Post_Data = 8'hC4; 
	12'hAB9 : Post_Data = 8'hC4; 
	12'hABA : Post_Data = 8'hC4; 
	12'hABB : Post_Data = 8'hC4; 
	12'hABC : Post_Data = 8'hC4; 
	12'hABD : Post_Data = 8'hC4; 
	12'hABE : Post_Data = 8'hC4; 
	12'hABF : Post_Data = 8'hC4; 
	12'hAC0 : Post_Data = 8'hC4; 
	12'hAC1 : Post_Data = 8'hC4; 
	12'hAC2 : Post_Data = 8'hC5; 
	12'hAC3 : Post_Data = 8'hC5; 
	12'hAC4 : Post_Data = 8'hC5; 
	12'hAC5 : Post_Data = 8'hC5; 
	12'hAC6 : Post_Data = 8'hC5; 
	12'hAC7 : Post_Data = 8'hC5; 
	12'hAC8 : Post_Data = 8'hC5; 
	12'hAC9 : Post_Data = 8'hC5; 
	12'hACA : Post_Data = 8'hC5; 
	12'hACB : Post_Data = 8'hC5; 
	12'hACC : Post_Data = 8'hC5; 
	12'hACD : Post_Data = 8'hC5; 
	12'hACE : Post_Data = 8'hC5; 
	12'hACF : Post_Data = 8'hC5; 
	12'hAD0 : Post_Data = 8'hC5; 
	12'hAD1 : Post_Data = 8'hC5; 
	12'hAD2 : Post_Data = 8'hC5; 
	12'hAD3 : Post_Data = 8'hC5; 
	12'hAD4 : Post_Data = 8'hC5; 
	12'hAD5 : Post_Data = 8'hC5; 
	12'hAD6 : Post_Data = 8'hC5; 
	12'hAD7 : Post_Data = 8'hC6; 
	12'hAD8 : Post_Data = 8'hC6; 
	12'hAD9 : Post_Data = 8'hC6; 
	12'hADA : Post_Data = 8'hC6; 
	12'hADB : Post_Data = 8'hC6; 
	12'hADC : Post_Data = 8'hC6; 
	12'hADD : Post_Data = 8'hC6; 
	12'hADE : Post_Data = 8'hC6; 
	12'hADF : Post_Data = 8'hC6; 
	12'hAE0 : Post_Data = 8'hC6; 
	12'hAE1 : Post_Data = 8'hC6; 
	12'hAE2 : Post_Data = 8'hC6; 
	12'hAE3 : Post_Data = 8'hC6; 
	12'hAE4 : Post_Data = 8'hC6; 
	12'hAE5 : Post_Data = 8'hC6; 
	12'hAE6 : Post_Data = 8'hC6; 
	12'hAE7 : Post_Data = 8'hC6; 
	12'hAE8 : Post_Data = 8'hC6; 
	12'hAE9 : Post_Data = 8'hC6; 
	12'hAEA : Post_Data = 8'hC6; 
	12'hAEB : Post_Data = 8'hC6; 
	12'hAEC : Post_Data = 8'hC7; 
	12'hAED : Post_Data = 8'hC7; 
	12'hAEE : Post_Data = 8'hC7; 
	12'hAEF : Post_Data = 8'hC7; 
	12'hAF0 : Post_Data = 8'hC7; 
	12'hAF1 : Post_Data = 8'hC7; 
	12'hAF2 : Post_Data = 8'hC7; 
	12'hAF3 : Post_Data = 8'hC7; 
	12'hAF4 : Post_Data = 8'hC7; 
	12'hAF5 : Post_Data = 8'hC7; 
	12'hAF6 : Post_Data = 8'hC7; 
	12'hAF7 : Post_Data = 8'hC7; 
	12'hAF8 : Post_Data = 8'hC7; 
	12'hAF9 : Post_Data = 8'hC7; 
	12'hAFA : Post_Data = 8'hC7; 
	12'hAFB : Post_Data = 8'hC7; 
	12'hAFC : Post_Data = 8'hC7; 
	12'hAFD : Post_Data = 8'hC7; 
	12'hAFE : Post_Data = 8'hC7; 
	12'hAFF : Post_Data = 8'hC7; 
	12'hB00 : Post_Data = 8'hC7; 
	12'hB01 : Post_Data = 8'hC8; 
	12'hB02 : Post_Data = 8'hC8; 
	12'hB03 : Post_Data = 8'hC8; 
	12'hB04 : Post_Data = 8'hC8; 
	12'hB05 : Post_Data = 8'hC8; 
	12'hB06 : Post_Data = 8'hC8; 
	12'hB07 : Post_Data = 8'hC8; 
	12'hB08 : Post_Data = 8'hC8; 
	12'hB09 : Post_Data = 8'hC8; 
	12'hB0A : Post_Data = 8'hC8; 
	12'hB0B : Post_Data = 8'hC8; 
	12'hB0C : Post_Data = 8'hC8; 
	12'hB0D : Post_Data = 8'hC8; 
	12'hB0E : Post_Data = 8'hC8; 
	12'hB0F : Post_Data = 8'hC8; 
	12'hB10 : Post_Data = 8'hC8; 
	12'hB11 : Post_Data = 8'hC8; 
	12'hB12 : Post_Data = 8'hC8; 
	12'hB13 : Post_Data = 8'hC8; 
	12'hB14 : Post_Data = 8'hC8; 
	12'hB15 : Post_Data = 8'hC8; 
	12'hB16 : Post_Data = 8'hC8; 
	12'hB17 : Post_Data = 8'hC9; 
	12'hB18 : Post_Data = 8'hC9; 
	12'hB19 : Post_Data = 8'hC9; 
	12'hB1A : Post_Data = 8'hC9; 
	12'hB1B : Post_Data = 8'hC9; 
	12'hB1C : Post_Data = 8'hC9; 
	12'hB1D : Post_Data = 8'hC9; 
	12'hB1E : Post_Data = 8'hC9; 
	12'hB1F : Post_Data = 8'hC9; 
	12'hB20 : Post_Data = 8'hC9; 
	12'hB21 : Post_Data = 8'hC9; 
	12'hB22 : Post_Data = 8'hC9; 
	12'hB23 : Post_Data = 8'hC9; 
	12'hB24 : Post_Data = 8'hC9; 
	12'hB25 : Post_Data = 8'hC9; 
	12'hB26 : Post_Data = 8'hC9; 
	12'hB27 : Post_Data = 8'hC9; 
	12'hB28 : Post_Data = 8'hC9; 
	12'hB29 : Post_Data = 8'hC9; 
	12'hB2A : Post_Data = 8'hC9; 
	12'hB2B : Post_Data = 8'hC9; 
	12'hB2C : Post_Data = 8'hCA; 
	12'hB2D : Post_Data = 8'hCA; 
	12'hB2E : Post_Data = 8'hCA; 
	12'hB2F : Post_Data = 8'hCA; 
	12'hB30 : Post_Data = 8'hCA; 
	12'hB31 : Post_Data = 8'hCA; 
	12'hB32 : Post_Data = 8'hCA; 
	12'hB33 : Post_Data = 8'hCA; 
	12'hB34 : Post_Data = 8'hCA; 
	12'hB35 : Post_Data = 8'hCA; 
	12'hB36 : Post_Data = 8'hCA; 
	12'hB37 : Post_Data = 8'hCA; 
	12'hB38 : Post_Data = 8'hCA; 
	12'hB39 : Post_Data = 8'hCA; 
	12'hB3A : Post_Data = 8'hCA; 
	12'hB3B : Post_Data = 8'hCA; 
	12'hB3C : Post_Data = 8'hCA; 
	12'hB3D : Post_Data = 8'hCA; 
	12'hB3E : Post_Data = 8'hCA; 
	12'hB3F : Post_Data = 8'hCA; 
	12'hB40 : Post_Data = 8'hCA; 
	12'hB41 : Post_Data = 8'hCB; 
	12'hB42 : Post_Data = 8'hCB; 
	12'hB43 : Post_Data = 8'hCB; 
	12'hB44 : Post_Data = 8'hCB; 
	12'hB45 : Post_Data = 8'hCB; 
	12'hB46 : Post_Data = 8'hCB; 
	12'hB47 : Post_Data = 8'hCB; 
	12'hB48 : Post_Data = 8'hCB; 
	12'hB49 : Post_Data = 8'hCB; 
	12'hB4A : Post_Data = 8'hCB; 
	12'hB4B : Post_Data = 8'hCB; 
	12'hB4C : Post_Data = 8'hCB; 
	12'hB4D : Post_Data = 8'hCB; 
	12'hB4E : Post_Data = 8'hCB; 
	12'hB4F : Post_Data = 8'hCB; 
	12'hB50 : Post_Data = 8'hCB; 
	12'hB51 : Post_Data = 8'hCB; 
	12'hB52 : Post_Data = 8'hCB; 
	12'hB53 : Post_Data = 8'hCB; 
	12'hB54 : Post_Data = 8'hCB; 
	12'hB55 : Post_Data = 8'hCB; 
	12'hB56 : Post_Data = 8'hCC; 
	12'hB57 : Post_Data = 8'hCC; 
	12'hB58 : Post_Data = 8'hCC; 
	12'hB59 : Post_Data = 8'hCC; 
	12'hB5A : Post_Data = 8'hCC; 
	12'hB5B : Post_Data = 8'hCC; 
	12'hB5C : Post_Data = 8'hCC; 
	12'hB5D : Post_Data = 8'hCC; 
	12'hB5E : Post_Data = 8'hCC; 
	12'hB5F : Post_Data = 8'hCC; 
	12'hB60 : Post_Data = 8'hCC; 
	12'hB61 : Post_Data = 8'hCC; 
	12'hB62 : Post_Data = 8'hCC; 
	12'hB63 : Post_Data = 8'hCC; 
	12'hB64 : Post_Data = 8'hCC; 
	12'hB65 : Post_Data = 8'hCC; 
	12'hB66 : Post_Data = 8'hCC; 
	12'hB67 : Post_Data = 8'hCC; 
	12'hB68 : Post_Data = 8'hCC; 
	12'hB69 : Post_Data = 8'hCC; 
	12'hB6A : Post_Data = 8'hCC; 
	12'hB6B : Post_Data = 8'hCC; 
	12'hB6C : Post_Data = 8'hCD; 
	12'hB6D : Post_Data = 8'hCD; 
	12'hB6E : Post_Data = 8'hCD; 
	12'hB6F : Post_Data = 8'hCD; 
	12'hB70 : Post_Data = 8'hCD; 
	12'hB71 : Post_Data = 8'hCD; 
	12'hB72 : Post_Data = 8'hCD; 
	12'hB73 : Post_Data = 8'hCD; 
	12'hB74 : Post_Data = 8'hCD; 
	12'hB75 : Post_Data = 8'hCD; 
	12'hB76 : Post_Data = 8'hCD; 
	12'hB77 : Post_Data = 8'hCD; 
	12'hB78 : Post_Data = 8'hCD; 
	12'hB79 : Post_Data = 8'hCD; 
	12'hB7A : Post_Data = 8'hCD; 
	12'hB7B : Post_Data = 8'hCD; 
	12'hB7C : Post_Data = 8'hCD; 
	12'hB7D : Post_Data = 8'hCD; 
	12'hB7E : Post_Data = 8'hCD; 
	12'hB7F : Post_Data = 8'hCD; 
	12'hB80 : Post_Data = 8'hCD; 
	12'hB81 : Post_Data = 8'hCE; 
	12'hB82 : Post_Data = 8'hCE; 
	12'hB83 : Post_Data = 8'hCE; 
	12'hB84 : Post_Data = 8'hCE; 
	12'hB85 : Post_Data = 8'hCE; 
	12'hB86 : Post_Data = 8'hCE; 
	12'hB87 : Post_Data = 8'hCE; 
	12'hB88 : Post_Data = 8'hCE; 
	12'hB89 : Post_Data = 8'hCE; 
	12'hB8A : Post_Data = 8'hCE; 
	12'hB8B : Post_Data = 8'hCE; 
	12'hB8C : Post_Data = 8'hCE; 
	12'hB8D : Post_Data = 8'hCE; 
	12'hB8E : Post_Data = 8'hCE; 
	12'hB8F : Post_Data = 8'hCE; 
	12'hB90 : Post_Data = 8'hCE; 
	12'hB91 : Post_Data = 8'hCE; 
	12'hB92 : Post_Data = 8'hCE; 
	12'hB93 : Post_Data = 8'hCE; 
	12'hB94 : Post_Data = 8'hCE; 
	12'hB95 : Post_Data = 8'hCE; 
	12'hB96 : Post_Data = 8'hCE; 
	12'hB97 : Post_Data = 8'hCF; 
	12'hB98 : Post_Data = 8'hCF; 
	12'hB99 : Post_Data = 8'hCF; 
	12'hB9A : Post_Data = 8'hCF; 
	12'hB9B : Post_Data = 8'hCF; 
	12'hB9C : Post_Data = 8'hCF; 
	12'hB9D : Post_Data = 8'hCF; 
	12'hB9E : Post_Data = 8'hCF; 
	12'hB9F : Post_Data = 8'hCF; 
	12'hBA0 : Post_Data = 8'hCF; 
	12'hBA1 : Post_Data = 8'hCF; 
	12'hBA2 : Post_Data = 8'hCF; 
	12'hBA3 : Post_Data = 8'hCF; 
	12'hBA4 : Post_Data = 8'hCF; 
	12'hBA5 : Post_Data = 8'hCF; 
	12'hBA6 : Post_Data = 8'hCF; 
	12'hBA7 : Post_Data = 8'hCF; 
	12'hBA8 : Post_Data = 8'hCF; 
	12'hBA9 : Post_Data = 8'hCF; 
	12'hBAA : Post_Data = 8'hCF; 
	12'hBAB : Post_Data = 8'hCF; 
	12'hBAC : Post_Data = 8'hCF; 
	12'hBAD : Post_Data = 8'hD0; 
	12'hBAE : Post_Data = 8'hD0; 
	12'hBAF : Post_Data = 8'hD0; 
	12'hBB0 : Post_Data = 8'hD0; 
	12'hBB1 : Post_Data = 8'hD0; 
	12'hBB2 : Post_Data = 8'hD0; 
	12'hBB3 : Post_Data = 8'hD0; 
	12'hBB4 : Post_Data = 8'hD0; 
	12'hBB5 : Post_Data = 8'hD0; 
	12'hBB6 : Post_Data = 8'hD0; 
	12'hBB7 : Post_Data = 8'hD0; 
	12'hBB8 : Post_Data = 8'hD0; 
	12'hBB9 : Post_Data = 8'hD0; 
	12'hBBA : Post_Data = 8'hD0; 
	12'hBBB : Post_Data = 8'hD0; 
	12'hBBC : Post_Data = 8'hD0; 
	12'hBBD : Post_Data = 8'hD0; 
	12'hBBE : Post_Data = 8'hD0; 
	12'hBBF : Post_Data = 8'hD0; 
	12'hBC0 : Post_Data = 8'hD0; 
	12'hBC1 : Post_Data = 8'hD0; 
	12'hBC2 : Post_Data = 8'hD1; 
	12'hBC3 : Post_Data = 8'hD1; 
	12'hBC4 : Post_Data = 8'hD1; 
	12'hBC5 : Post_Data = 8'hD1; 
	12'hBC6 : Post_Data = 8'hD1; 
	12'hBC7 : Post_Data = 8'hD1; 
	12'hBC8 : Post_Data = 8'hD1; 
	12'hBC9 : Post_Data = 8'hD1; 
	12'hBCA : Post_Data = 8'hD1; 
	12'hBCB : Post_Data = 8'hD1; 
	12'hBCC : Post_Data = 8'hD1; 
	12'hBCD : Post_Data = 8'hD1; 
	12'hBCE : Post_Data = 8'hD1; 
	12'hBCF : Post_Data = 8'hD1; 
	12'hBD0 : Post_Data = 8'hD1; 
	12'hBD1 : Post_Data = 8'hD1; 
	12'hBD2 : Post_Data = 8'hD1; 
	12'hBD3 : Post_Data = 8'hD1; 
	12'hBD4 : Post_Data = 8'hD1; 
	12'hBD5 : Post_Data = 8'hD1; 
	12'hBD6 : Post_Data = 8'hD1; 
	12'hBD7 : Post_Data = 8'hD1; 
	12'hBD8 : Post_Data = 8'hD2; 
	12'hBD9 : Post_Data = 8'hD2; 
	12'hBDA : Post_Data = 8'hD2; 
	12'hBDB : Post_Data = 8'hD2; 
	12'hBDC : Post_Data = 8'hD2; 
	12'hBDD : Post_Data = 8'hD2; 
	12'hBDE : Post_Data = 8'hD2; 
	12'hBDF : Post_Data = 8'hD2; 
	12'hBE0 : Post_Data = 8'hD2; 
	12'hBE1 : Post_Data = 8'hD2; 
	12'hBE2 : Post_Data = 8'hD2; 
	12'hBE3 : Post_Data = 8'hD2; 
	12'hBE4 : Post_Data = 8'hD2; 
	12'hBE5 : Post_Data = 8'hD2; 
	12'hBE6 : Post_Data = 8'hD2; 
	12'hBE7 : Post_Data = 8'hD2; 
	12'hBE8 : Post_Data = 8'hD2; 
	12'hBE9 : Post_Data = 8'hD2; 
	12'hBEA : Post_Data = 8'hD2; 
	12'hBEB : Post_Data = 8'hD2; 
	12'hBEC : Post_Data = 8'hD2; 
	12'hBED : Post_Data = 8'hD2; 
	12'hBEE : Post_Data = 8'hD3; 
	12'hBEF : Post_Data = 8'hD3; 
	12'hBF0 : Post_Data = 8'hD3; 
	12'hBF1 : Post_Data = 8'hD3; 
	12'hBF2 : Post_Data = 8'hD3; 
	12'hBF3 : Post_Data = 8'hD3; 
	12'hBF4 : Post_Data = 8'hD3; 
	12'hBF5 : Post_Data = 8'hD3; 
	12'hBF6 : Post_Data = 8'hD3; 
	12'hBF7 : Post_Data = 8'hD3; 
	12'hBF8 : Post_Data = 8'hD3; 
	12'hBF9 : Post_Data = 8'hD3; 
	12'hBFA : Post_Data = 8'hD3; 
	12'hBFB : Post_Data = 8'hD3; 
	12'hBFC : Post_Data = 8'hD3; 
	12'hBFD : Post_Data = 8'hD3; 
	12'hBFE : Post_Data = 8'hD3; 
	12'hBFF : Post_Data = 8'hD3; 
	12'hC00 : Post_Data = 8'hD3; 
	12'hC01 : Post_Data = 8'hD3; 
	12'hC02 : Post_Data = 8'hD3; 
	12'hC03 : Post_Data = 8'hD4; 
	12'hC04 : Post_Data = 8'hD4; 
	12'hC05 : Post_Data = 8'hD4; 
	12'hC06 : Post_Data = 8'hD4; 
	12'hC07 : Post_Data = 8'hD4; 
	12'hC08 : Post_Data = 8'hD4; 
	12'hC09 : Post_Data = 8'hD4; 
	12'hC0A : Post_Data = 8'hD4; 
	12'hC0B : Post_Data = 8'hD4; 
	12'hC0C : Post_Data = 8'hD4; 
	12'hC0D : Post_Data = 8'hD4; 
	12'hC0E : Post_Data = 8'hD4; 
	12'hC0F : Post_Data = 8'hD4; 
	12'hC10 : Post_Data = 8'hD4; 
	12'hC11 : Post_Data = 8'hD4; 
	12'hC12 : Post_Data = 8'hD4; 
	12'hC13 : Post_Data = 8'hD4; 
	12'hC14 : Post_Data = 8'hD4; 
	12'hC15 : Post_Data = 8'hD4; 
	12'hC16 : Post_Data = 8'hD4; 
	12'hC17 : Post_Data = 8'hD4; 
	12'hC18 : Post_Data = 8'hD4; 
	12'hC19 : Post_Data = 8'hD5; 
	12'hC1A : Post_Data = 8'hD5; 
	12'hC1B : Post_Data = 8'hD5; 
	12'hC1C : Post_Data = 8'hD5; 
	12'hC1D : Post_Data = 8'hD5; 
	12'hC1E : Post_Data = 8'hD5; 
	12'hC1F : Post_Data = 8'hD5; 
	12'hC20 : Post_Data = 8'hD5; 
	12'hC21 : Post_Data = 8'hD5; 
	12'hC22 : Post_Data = 8'hD5; 
	12'hC23 : Post_Data = 8'hD5; 
	12'hC24 : Post_Data = 8'hD5; 
	12'hC25 : Post_Data = 8'hD5; 
	12'hC26 : Post_Data = 8'hD5; 
	12'hC27 : Post_Data = 8'hD5; 
	12'hC28 : Post_Data = 8'hD5; 
	12'hC29 : Post_Data = 8'hD5; 
	12'hC2A : Post_Data = 8'hD5; 
	12'hC2B : Post_Data = 8'hD5; 
	12'hC2C : Post_Data = 8'hD5; 
	12'hC2D : Post_Data = 8'hD5; 
	12'hC2E : Post_Data = 8'hD5; 
	12'hC2F : Post_Data = 8'hD6; 
	12'hC30 : Post_Data = 8'hD6; 
	12'hC31 : Post_Data = 8'hD6; 
	12'hC32 : Post_Data = 8'hD6; 
	12'hC33 : Post_Data = 8'hD6; 
	12'hC34 : Post_Data = 8'hD6; 
	12'hC35 : Post_Data = 8'hD6; 
	12'hC36 : Post_Data = 8'hD6; 
	12'hC37 : Post_Data = 8'hD6; 
	12'hC38 : Post_Data = 8'hD6; 
	12'hC39 : Post_Data = 8'hD6; 
	12'hC3A : Post_Data = 8'hD6; 
	12'hC3B : Post_Data = 8'hD6; 
	12'hC3C : Post_Data = 8'hD6; 
	12'hC3D : Post_Data = 8'hD6; 
	12'hC3E : Post_Data = 8'hD6; 
	12'hC3F : Post_Data = 8'hD6; 
	12'hC40 : Post_Data = 8'hD6; 
	12'hC41 : Post_Data = 8'hD6; 
	12'hC42 : Post_Data = 8'hD6; 
	12'hC43 : Post_Data = 8'hD6; 
	12'hC44 : Post_Data = 8'hD6; 
	12'hC45 : Post_Data = 8'hD7; 
	12'hC46 : Post_Data = 8'hD7; 
	12'hC47 : Post_Data = 8'hD7; 
	12'hC48 : Post_Data = 8'hD7; 
	12'hC49 : Post_Data = 8'hD7; 
	12'hC4A : Post_Data = 8'hD7; 
	12'hC4B : Post_Data = 8'hD7; 
	12'hC4C : Post_Data = 8'hD7; 
	12'hC4D : Post_Data = 8'hD7; 
	12'hC4E : Post_Data = 8'hD7; 
	12'hC4F : Post_Data = 8'hD7; 
	12'hC50 : Post_Data = 8'hD7; 
	12'hC51 : Post_Data = 8'hD7; 
	12'hC52 : Post_Data = 8'hD7; 
	12'hC53 : Post_Data = 8'hD7; 
	12'hC54 : Post_Data = 8'hD7; 
	12'hC55 : Post_Data = 8'hD7; 
	12'hC56 : Post_Data = 8'hD7; 
	12'hC57 : Post_Data = 8'hD7; 
	12'hC58 : Post_Data = 8'hD7; 
	12'hC59 : Post_Data = 8'hD7; 
	12'hC5A : Post_Data = 8'hD7; 
	12'hC5B : Post_Data = 8'hD8; 
	12'hC5C : Post_Data = 8'hD8; 
	12'hC5D : Post_Data = 8'hD8; 
	12'hC5E : Post_Data = 8'hD8; 
	12'hC5F : Post_Data = 8'hD8; 
	12'hC60 : Post_Data = 8'hD8; 
	12'hC61 : Post_Data = 8'hD8; 
	12'hC62 : Post_Data = 8'hD8; 
	12'hC63 : Post_Data = 8'hD8; 
	12'hC64 : Post_Data = 8'hD8; 
	12'hC65 : Post_Data = 8'hD8; 
	12'hC66 : Post_Data = 8'hD8; 
	12'hC67 : Post_Data = 8'hD8; 
	12'hC68 : Post_Data = 8'hD8; 
	12'hC69 : Post_Data = 8'hD8; 
	12'hC6A : Post_Data = 8'hD8; 
	12'hC6B : Post_Data = 8'hD8; 
	12'hC6C : Post_Data = 8'hD8; 
	12'hC6D : Post_Data = 8'hD8; 
	12'hC6E : Post_Data = 8'hD8; 
	12'hC6F : Post_Data = 8'hD8; 
	12'hC70 : Post_Data = 8'hD8; 
	12'hC71 : Post_Data = 8'hD9; 
	12'hC72 : Post_Data = 8'hD9; 
	12'hC73 : Post_Data = 8'hD9; 
	12'hC74 : Post_Data = 8'hD9; 
	12'hC75 : Post_Data = 8'hD9; 
	12'hC76 : Post_Data = 8'hD9; 
	12'hC77 : Post_Data = 8'hD9; 
	12'hC78 : Post_Data = 8'hD9; 
	12'hC79 : Post_Data = 8'hD9; 
	12'hC7A : Post_Data = 8'hD9; 
	12'hC7B : Post_Data = 8'hD9; 
	12'hC7C : Post_Data = 8'hD9; 
	12'hC7D : Post_Data = 8'hD9; 
	12'hC7E : Post_Data = 8'hD9; 
	12'hC7F : Post_Data = 8'hD9; 
	12'hC80 : Post_Data = 8'hD9; 
	12'hC81 : Post_Data = 8'hD9; 
	12'hC82 : Post_Data = 8'hD9; 
	12'hC83 : Post_Data = 8'hD9; 
	12'hC84 : Post_Data = 8'hD9; 
	12'hC85 : Post_Data = 8'hD9; 
	12'hC86 : Post_Data = 8'hD9; 
	12'hC87 : Post_Data = 8'hDA; 
	12'hC88 : Post_Data = 8'hDA; 
	12'hC89 : Post_Data = 8'hDA; 
	12'hC8A : Post_Data = 8'hDA; 
	12'hC8B : Post_Data = 8'hDA; 
	12'hC8C : Post_Data = 8'hDA; 
	12'hC8D : Post_Data = 8'hDA; 
	12'hC8E : Post_Data = 8'hDA; 
	12'hC8F : Post_Data = 8'hDA; 
	12'hC90 : Post_Data = 8'hDA; 
	12'hC91 : Post_Data = 8'hDA; 
	12'hC92 : Post_Data = 8'hDA; 
	12'hC93 : Post_Data = 8'hDA; 
	12'hC94 : Post_Data = 8'hDA; 
	12'hC95 : Post_Data = 8'hDA; 
	12'hC96 : Post_Data = 8'hDA; 
	12'hC97 : Post_Data = 8'hDA; 
	12'hC98 : Post_Data = 8'hDA; 
	12'hC99 : Post_Data = 8'hDA; 
	12'hC9A : Post_Data = 8'hDA; 
	12'hC9B : Post_Data = 8'hDA; 
	12'hC9C : Post_Data = 8'hDA; 
	12'hC9D : Post_Data = 8'hDB; 
	12'hC9E : Post_Data = 8'hDB; 
	12'hC9F : Post_Data = 8'hDB; 
	12'hCA0 : Post_Data = 8'hDB; 
	12'hCA1 : Post_Data = 8'hDB; 
	12'hCA2 : Post_Data = 8'hDB; 
	12'hCA3 : Post_Data = 8'hDB; 
	12'hCA4 : Post_Data = 8'hDB; 
	12'hCA5 : Post_Data = 8'hDB; 
	12'hCA6 : Post_Data = 8'hDB; 
	12'hCA7 : Post_Data = 8'hDB; 
	12'hCA8 : Post_Data = 8'hDB; 
	12'hCA9 : Post_Data = 8'hDB; 
	12'hCAA : Post_Data = 8'hDB; 
	12'hCAB : Post_Data = 8'hDB; 
	12'hCAC : Post_Data = 8'hDB; 
	12'hCAD : Post_Data = 8'hDB; 
	12'hCAE : Post_Data = 8'hDB; 
	12'hCAF : Post_Data = 8'hDB; 
	12'hCB0 : Post_Data = 8'hDB; 
	12'hCB1 : Post_Data = 8'hDB; 
	12'hCB2 : Post_Data = 8'hDB; 
	12'hCB3 : Post_Data = 8'hDB; 
	12'hCB4 : Post_Data = 8'hDC; 
	12'hCB5 : Post_Data = 8'hDC; 
	12'hCB6 : Post_Data = 8'hDC; 
	12'hCB7 : Post_Data = 8'hDC; 
	12'hCB8 : Post_Data = 8'hDC; 
	12'hCB9 : Post_Data = 8'hDC; 
	12'hCBA : Post_Data = 8'hDC; 
	12'hCBB : Post_Data = 8'hDC; 
	12'hCBC : Post_Data = 8'hDC; 
	12'hCBD : Post_Data = 8'hDC; 
	12'hCBE : Post_Data = 8'hDC; 
	12'hCBF : Post_Data = 8'hDC; 
	12'hCC0 : Post_Data = 8'hDC; 
	12'hCC1 : Post_Data = 8'hDC; 
	12'hCC2 : Post_Data = 8'hDC; 
	12'hCC3 : Post_Data = 8'hDC; 
	12'hCC4 : Post_Data = 8'hDC; 
	12'hCC5 : Post_Data = 8'hDC; 
	12'hCC6 : Post_Data = 8'hDC; 
	12'hCC7 : Post_Data = 8'hDC; 
	12'hCC8 : Post_Data = 8'hDC; 
	12'hCC9 : Post_Data = 8'hDC; 
	12'hCCA : Post_Data = 8'hDD; 
	12'hCCB : Post_Data = 8'hDD; 
	12'hCCC : Post_Data = 8'hDD; 
	12'hCCD : Post_Data = 8'hDD; 
	12'hCCE : Post_Data = 8'hDD; 
	12'hCCF : Post_Data = 8'hDD; 
	12'hCD0 : Post_Data = 8'hDD; 
	12'hCD1 : Post_Data = 8'hDD; 
	12'hCD2 : Post_Data = 8'hDD; 
	12'hCD3 : Post_Data = 8'hDD; 
	12'hCD4 : Post_Data = 8'hDD; 
	12'hCD5 : Post_Data = 8'hDD; 
	12'hCD6 : Post_Data = 8'hDD; 
	12'hCD7 : Post_Data = 8'hDD; 
	12'hCD8 : Post_Data = 8'hDD; 
	12'hCD9 : Post_Data = 8'hDD; 
	12'hCDA : Post_Data = 8'hDD; 
	12'hCDB : Post_Data = 8'hDD; 
	12'hCDC : Post_Data = 8'hDD; 
	12'hCDD : Post_Data = 8'hDD; 
	12'hCDE : Post_Data = 8'hDD; 
	12'hCDF : Post_Data = 8'hDD; 
	12'hCE0 : Post_Data = 8'hDE; 
	12'hCE1 : Post_Data = 8'hDE; 
	12'hCE2 : Post_Data = 8'hDE; 
	12'hCE3 : Post_Data = 8'hDE; 
	12'hCE4 : Post_Data = 8'hDE; 
	12'hCE5 : Post_Data = 8'hDE; 
	12'hCE6 : Post_Data = 8'hDE; 
	12'hCE7 : Post_Data = 8'hDE; 
	12'hCE8 : Post_Data = 8'hDE; 
	12'hCE9 : Post_Data = 8'hDE; 
	12'hCEA : Post_Data = 8'hDE; 
	12'hCEB : Post_Data = 8'hDE; 
	12'hCEC : Post_Data = 8'hDE; 
	12'hCED : Post_Data = 8'hDE; 
	12'hCEE : Post_Data = 8'hDE; 
	12'hCEF : Post_Data = 8'hDE; 
	12'hCF0 : Post_Data = 8'hDE; 
	12'hCF1 : Post_Data = 8'hDE; 
	12'hCF2 : Post_Data = 8'hDE; 
	12'hCF3 : Post_Data = 8'hDE; 
	12'hCF4 : Post_Data = 8'hDE; 
	12'hCF5 : Post_Data = 8'hDE; 
	12'hCF6 : Post_Data = 8'hDF; 
	12'hCF7 : Post_Data = 8'hDF; 
	12'hCF8 : Post_Data = 8'hDF; 
	12'hCF9 : Post_Data = 8'hDF; 
	12'hCFA : Post_Data = 8'hDF; 
	12'hCFB : Post_Data = 8'hDF; 
	12'hCFC : Post_Data = 8'hDF; 
	12'hCFD : Post_Data = 8'hDF; 
	12'hCFE : Post_Data = 8'hDF; 
	12'hCFF : Post_Data = 8'hDF; 
	12'hD00 : Post_Data = 8'hDF; 
	12'hD01 : Post_Data = 8'hDF; 
	12'hD02 : Post_Data = 8'hDF; 
	12'hD03 : Post_Data = 8'hDF; 
	12'hD04 : Post_Data = 8'hDF; 
	12'hD05 : Post_Data = 8'hDF; 
	12'hD06 : Post_Data = 8'hDF; 
	12'hD07 : Post_Data = 8'hDF; 
	12'hD08 : Post_Data = 8'hDF; 
	12'hD09 : Post_Data = 8'hDF; 
	12'hD0A : Post_Data = 8'hDF; 
	12'hD0B : Post_Data = 8'hDF; 
	12'hD0C : Post_Data = 8'hDF; 
	12'hD0D : Post_Data = 8'hE0; 
	12'hD0E : Post_Data = 8'hE0; 
	12'hD0F : Post_Data = 8'hE0; 
	12'hD10 : Post_Data = 8'hE0; 
	12'hD11 : Post_Data = 8'hE0; 
	12'hD12 : Post_Data = 8'hE0; 
	12'hD13 : Post_Data = 8'hE0; 
	12'hD14 : Post_Data = 8'hE0; 
	12'hD15 : Post_Data = 8'hE0; 
	12'hD16 : Post_Data = 8'hE0; 
	12'hD17 : Post_Data = 8'hE0; 
	12'hD18 : Post_Data = 8'hE0; 
	12'hD19 : Post_Data = 8'hE0; 
	12'hD1A : Post_Data = 8'hE0; 
	12'hD1B : Post_Data = 8'hE0; 
	12'hD1C : Post_Data = 8'hE0; 
	12'hD1D : Post_Data = 8'hE0; 
	12'hD1E : Post_Data = 8'hE0; 
	12'hD1F : Post_Data = 8'hE0; 
	12'hD20 : Post_Data = 8'hE0; 
	12'hD21 : Post_Data = 8'hE0; 
	12'hD22 : Post_Data = 8'hE0; 
	12'hD23 : Post_Data = 8'hE1; 
	12'hD24 : Post_Data = 8'hE1; 
	12'hD25 : Post_Data = 8'hE1; 
	12'hD26 : Post_Data = 8'hE1; 
	12'hD27 : Post_Data = 8'hE1; 
	12'hD28 : Post_Data = 8'hE1; 
	12'hD29 : Post_Data = 8'hE1; 
	12'hD2A : Post_Data = 8'hE1; 
	12'hD2B : Post_Data = 8'hE1; 
	12'hD2C : Post_Data = 8'hE1; 
	12'hD2D : Post_Data = 8'hE1; 
	12'hD2E : Post_Data = 8'hE1; 
	12'hD2F : Post_Data = 8'hE1; 
	12'hD30 : Post_Data = 8'hE1; 
	12'hD31 : Post_Data = 8'hE1; 
	12'hD32 : Post_Data = 8'hE1; 
	12'hD33 : Post_Data = 8'hE1; 
	12'hD34 : Post_Data = 8'hE1; 
	12'hD35 : Post_Data = 8'hE1; 
	12'hD36 : Post_Data = 8'hE1; 
	12'hD37 : Post_Data = 8'hE1; 
	12'hD38 : Post_Data = 8'hE1; 
	12'hD39 : Post_Data = 8'hE1; 
	12'hD3A : Post_Data = 8'hE2; 
	12'hD3B : Post_Data = 8'hE2; 
	12'hD3C : Post_Data = 8'hE2; 
	12'hD3D : Post_Data = 8'hE2; 
	12'hD3E : Post_Data = 8'hE2; 
	12'hD3F : Post_Data = 8'hE2; 
	12'hD40 : Post_Data = 8'hE2; 
	12'hD41 : Post_Data = 8'hE2; 
	12'hD42 : Post_Data = 8'hE2; 
	12'hD43 : Post_Data = 8'hE2; 
	12'hD44 : Post_Data = 8'hE2; 
	12'hD45 : Post_Data = 8'hE2; 
	12'hD46 : Post_Data = 8'hE2; 
	12'hD47 : Post_Data = 8'hE2; 
	12'hD48 : Post_Data = 8'hE2; 
	12'hD49 : Post_Data = 8'hE2; 
	12'hD4A : Post_Data = 8'hE2; 
	12'hD4B : Post_Data = 8'hE2; 
	12'hD4C : Post_Data = 8'hE2; 
	12'hD4D : Post_Data = 8'hE2; 
	12'hD4E : Post_Data = 8'hE2; 
	12'hD4F : Post_Data = 8'hE2; 
	12'hD50 : Post_Data = 8'hE3; 
	12'hD51 : Post_Data = 8'hE3; 
	12'hD52 : Post_Data = 8'hE3; 
	12'hD53 : Post_Data = 8'hE3; 
	12'hD54 : Post_Data = 8'hE3; 
	12'hD55 : Post_Data = 8'hE3; 
	12'hD56 : Post_Data = 8'hE3; 
	12'hD57 : Post_Data = 8'hE3; 
	12'hD58 : Post_Data = 8'hE3; 
	12'hD59 : Post_Data = 8'hE3; 
	12'hD5A : Post_Data = 8'hE3; 
	12'hD5B : Post_Data = 8'hE3; 
	12'hD5C : Post_Data = 8'hE3; 
	12'hD5D : Post_Data = 8'hE3; 
	12'hD5E : Post_Data = 8'hE3; 
	12'hD5F : Post_Data = 8'hE3; 
	12'hD60 : Post_Data = 8'hE3; 
	12'hD61 : Post_Data = 8'hE3; 
	12'hD62 : Post_Data = 8'hE3; 
	12'hD63 : Post_Data = 8'hE3; 
	12'hD64 : Post_Data = 8'hE3; 
	12'hD65 : Post_Data = 8'hE3; 
	12'hD66 : Post_Data = 8'hE3; 
	12'hD67 : Post_Data = 8'hE4; 
	12'hD68 : Post_Data = 8'hE4; 
	12'hD69 : Post_Data = 8'hE4; 
	12'hD6A : Post_Data = 8'hE4; 
	12'hD6B : Post_Data = 8'hE4; 
	12'hD6C : Post_Data = 8'hE4; 
	12'hD6D : Post_Data = 8'hE4; 
	12'hD6E : Post_Data = 8'hE4; 
	12'hD6F : Post_Data = 8'hE4; 
	12'hD70 : Post_Data = 8'hE4; 
	12'hD71 : Post_Data = 8'hE4; 
	12'hD72 : Post_Data = 8'hE4; 
	12'hD73 : Post_Data = 8'hE4; 
	12'hD74 : Post_Data = 8'hE4; 
	12'hD75 : Post_Data = 8'hE4; 
	12'hD76 : Post_Data = 8'hE4; 
	12'hD77 : Post_Data = 8'hE4; 
	12'hD78 : Post_Data = 8'hE4; 
	12'hD79 : Post_Data = 8'hE4; 
	12'hD7A : Post_Data = 8'hE4; 
	12'hD7B : Post_Data = 8'hE4; 
	12'hD7C : Post_Data = 8'hE4; 
	12'hD7D : Post_Data = 8'hE4; 
	12'hD7E : Post_Data = 8'hE5; 
	12'hD7F : Post_Data = 8'hE5; 
	12'hD80 : Post_Data = 8'hE5; 
	12'hD81 : Post_Data = 8'hE5; 
	12'hD82 : Post_Data = 8'hE5; 
	12'hD83 : Post_Data = 8'hE5; 
	12'hD84 : Post_Data = 8'hE5; 
	12'hD85 : Post_Data = 8'hE5; 
	12'hD86 : Post_Data = 8'hE5; 
	12'hD87 : Post_Data = 8'hE5; 
	12'hD88 : Post_Data = 8'hE5; 
	12'hD89 : Post_Data = 8'hE5; 
	12'hD8A : Post_Data = 8'hE5; 
	12'hD8B : Post_Data = 8'hE5; 
	12'hD8C : Post_Data = 8'hE5; 
	12'hD8D : Post_Data = 8'hE5; 
	12'hD8E : Post_Data = 8'hE5; 
	12'hD8F : Post_Data = 8'hE5; 
	12'hD90 : Post_Data = 8'hE5; 
	12'hD91 : Post_Data = 8'hE5; 
	12'hD92 : Post_Data = 8'hE5; 
	12'hD93 : Post_Data = 8'hE5; 
	12'hD94 : Post_Data = 8'hE6; 
	12'hD95 : Post_Data = 8'hE6; 
	12'hD96 : Post_Data = 8'hE6; 
	12'hD97 : Post_Data = 8'hE6; 
	12'hD98 : Post_Data = 8'hE6; 
	12'hD99 : Post_Data = 8'hE6; 
	12'hD9A : Post_Data = 8'hE6; 
	12'hD9B : Post_Data = 8'hE6; 
	12'hD9C : Post_Data = 8'hE6; 
	12'hD9D : Post_Data = 8'hE6; 
	12'hD9E : Post_Data = 8'hE6; 
	12'hD9F : Post_Data = 8'hE6; 
	12'hDA0 : Post_Data = 8'hE6; 
	12'hDA1 : Post_Data = 8'hE6; 
	12'hDA2 : Post_Data = 8'hE6; 
	12'hDA3 : Post_Data = 8'hE6; 
	12'hDA4 : Post_Data = 8'hE6; 
	12'hDA5 : Post_Data = 8'hE6; 
	12'hDA6 : Post_Data = 8'hE6; 
	12'hDA7 : Post_Data = 8'hE6; 
	12'hDA8 : Post_Data = 8'hE6; 
	12'hDA9 : Post_Data = 8'hE6; 
	12'hDAA : Post_Data = 8'hE6; 
	12'hDAB : Post_Data = 8'hE7; 
	12'hDAC : Post_Data = 8'hE7; 
	12'hDAD : Post_Data = 8'hE7; 
	12'hDAE : Post_Data = 8'hE7; 
	12'hDAF : Post_Data = 8'hE7; 
	12'hDB0 : Post_Data = 8'hE7; 
	12'hDB1 : Post_Data = 8'hE7; 
	12'hDB2 : Post_Data = 8'hE7; 
	12'hDB3 : Post_Data = 8'hE7; 
	12'hDB4 : Post_Data = 8'hE7; 
	12'hDB5 : Post_Data = 8'hE7; 
	12'hDB6 : Post_Data = 8'hE7; 
	12'hDB7 : Post_Data = 8'hE7; 
	12'hDB8 : Post_Data = 8'hE7; 
	12'hDB9 : Post_Data = 8'hE7; 
	12'hDBA : Post_Data = 8'hE7; 
	12'hDBB : Post_Data = 8'hE7; 
	12'hDBC : Post_Data = 8'hE7; 
	12'hDBD : Post_Data = 8'hE7; 
	12'hDBE : Post_Data = 8'hE7; 
	12'hDBF : Post_Data = 8'hE7; 
	12'hDC0 : Post_Data = 8'hE7; 
	12'hDC1 : Post_Data = 8'hE7; 
	12'hDC2 : Post_Data = 8'hE8; 
	12'hDC3 : Post_Data = 8'hE8; 
	12'hDC4 : Post_Data = 8'hE8; 
	12'hDC5 : Post_Data = 8'hE8; 
	12'hDC6 : Post_Data = 8'hE8; 
	12'hDC7 : Post_Data = 8'hE8; 
	12'hDC8 : Post_Data = 8'hE8; 
	12'hDC9 : Post_Data = 8'hE8; 
	12'hDCA : Post_Data = 8'hE8; 
	12'hDCB : Post_Data = 8'hE8; 
	12'hDCC : Post_Data = 8'hE8; 
	12'hDCD : Post_Data = 8'hE8; 
	12'hDCE : Post_Data = 8'hE8; 
	12'hDCF : Post_Data = 8'hE8; 
	12'hDD0 : Post_Data = 8'hE8; 
	12'hDD1 : Post_Data = 8'hE8; 
	12'hDD2 : Post_Data = 8'hE8; 
	12'hDD3 : Post_Data = 8'hE8; 
	12'hDD4 : Post_Data = 8'hE8; 
	12'hDD5 : Post_Data = 8'hE8; 
	12'hDD6 : Post_Data = 8'hE8; 
	12'hDD7 : Post_Data = 8'hE8; 
	12'hDD8 : Post_Data = 8'hE8; 
	12'hDD9 : Post_Data = 8'hE9; 
	12'hDDA : Post_Data = 8'hE9; 
	12'hDDB : Post_Data = 8'hE9; 
	12'hDDC : Post_Data = 8'hE9; 
	12'hDDD : Post_Data = 8'hE9; 
	12'hDDE : Post_Data = 8'hE9; 
	12'hDDF : Post_Data = 8'hE9; 
	12'hDE0 : Post_Data = 8'hE9; 
	12'hDE1 : Post_Data = 8'hE9; 
	12'hDE2 : Post_Data = 8'hE9; 
	12'hDE3 : Post_Data = 8'hE9; 
	12'hDE4 : Post_Data = 8'hE9; 
	12'hDE5 : Post_Data = 8'hE9; 
	12'hDE6 : Post_Data = 8'hE9; 
	12'hDE7 : Post_Data = 8'hE9; 
	12'hDE8 : Post_Data = 8'hE9; 
	12'hDE9 : Post_Data = 8'hE9; 
	12'hDEA : Post_Data = 8'hE9; 
	12'hDEB : Post_Data = 8'hE9; 
	12'hDEC : Post_Data = 8'hE9; 
	12'hDED : Post_Data = 8'hE9; 
	12'hDEE : Post_Data = 8'hE9; 
	12'hDEF : Post_Data = 8'hE9; 
	12'hDF0 : Post_Data = 8'hEA; 
	12'hDF1 : Post_Data = 8'hEA; 
	12'hDF2 : Post_Data = 8'hEA; 
	12'hDF3 : Post_Data = 8'hEA; 
	12'hDF4 : Post_Data = 8'hEA; 
	12'hDF5 : Post_Data = 8'hEA; 
	12'hDF6 : Post_Data = 8'hEA; 
	12'hDF7 : Post_Data = 8'hEA; 
	12'hDF8 : Post_Data = 8'hEA; 
	12'hDF9 : Post_Data = 8'hEA; 
	12'hDFA : Post_Data = 8'hEA; 
	12'hDFB : Post_Data = 8'hEA; 
	12'hDFC : Post_Data = 8'hEA; 
	12'hDFD : Post_Data = 8'hEA; 
	12'hDFE : Post_Data = 8'hEA; 
	12'hDFF : Post_Data = 8'hEA; 
	12'hE00 : Post_Data = 8'hEA; 
	12'hE01 : Post_Data = 8'hEA; 
	12'hE02 : Post_Data = 8'hEA; 
	12'hE03 : Post_Data = 8'hEA; 
	12'hE04 : Post_Data = 8'hEA; 
	12'hE05 : Post_Data = 8'hEA; 
	12'hE06 : Post_Data = 8'hEB; 
	12'hE07 : Post_Data = 8'hEB; 
	12'hE08 : Post_Data = 8'hEB; 
	12'hE09 : Post_Data = 8'hEB; 
	12'hE0A : Post_Data = 8'hEB; 
	12'hE0B : Post_Data = 8'hEB; 
	12'hE0C : Post_Data = 8'hEB; 
	12'hE0D : Post_Data = 8'hEB; 
	12'hE0E : Post_Data = 8'hEB; 
	12'hE0F : Post_Data = 8'hEB; 
	12'hE10 : Post_Data = 8'hEB; 
	12'hE11 : Post_Data = 8'hEB; 
	12'hE12 : Post_Data = 8'hEB; 
	12'hE13 : Post_Data = 8'hEB; 
	12'hE14 : Post_Data = 8'hEB; 
	12'hE15 : Post_Data = 8'hEB; 
	12'hE16 : Post_Data = 8'hEB; 
	12'hE17 : Post_Data = 8'hEB; 
	12'hE18 : Post_Data = 8'hEB; 
	12'hE19 : Post_Data = 8'hEB; 
	12'hE1A : Post_Data = 8'hEB; 
	12'hE1B : Post_Data = 8'hEB; 
	12'hE1C : Post_Data = 8'hEB; 
	12'hE1D : Post_Data = 8'hEC; 
	12'hE1E : Post_Data = 8'hEC; 
	12'hE1F : Post_Data = 8'hEC; 
	12'hE20 : Post_Data = 8'hEC; 
	12'hE21 : Post_Data = 8'hEC; 
	12'hE22 : Post_Data = 8'hEC; 
	12'hE23 : Post_Data = 8'hEC; 
	12'hE24 : Post_Data = 8'hEC; 
	12'hE25 : Post_Data = 8'hEC; 
	12'hE26 : Post_Data = 8'hEC; 
	12'hE27 : Post_Data = 8'hEC; 
	12'hE28 : Post_Data = 8'hEC; 
	12'hE29 : Post_Data = 8'hEC; 
	12'hE2A : Post_Data = 8'hEC; 
	12'hE2B : Post_Data = 8'hEC; 
	12'hE2C : Post_Data = 8'hEC; 
	12'hE2D : Post_Data = 8'hEC; 
	12'hE2E : Post_Data = 8'hEC; 
	12'hE2F : Post_Data = 8'hEC; 
	12'hE30 : Post_Data = 8'hEC; 
	12'hE31 : Post_Data = 8'hEC; 
	12'hE32 : Post_Data = 8'hEC; 
	12'hE33 : Post_Data = 8'hEC; 
	12'hE34 : Post_Data = 8'hEC; 
	12'hE35 : Post_Data = 8'hED; 
	12'hE36 : Post_Data = 8'hED; 
	12'hE37 : Post_Data = 8'hED; 
	12'hE38 : Post_Data = 8'hED; 
	12'hE39 : Post_Data = 8'hED; 
	12'hE3A : Post_Data = 8'hED; 
	12'hE3B : Post_Data = 8'hED; 
	12'hE3C : Post_Data = 8'hED; 
	12'hE3D : Post_Data = 8'hED; 
	12'hE3E : Post_Data = 8'hED; 
	12'hE3F : Post_Data = 8'hED; 
	12'hE40 : Post_Data = 8'hED; 
	12'hE41 : Post_Data = 8'hED; 
	12'hE42 : Post_Data = 8'hED; 
	12'hE43 : Post_Data = 8'hED; 
	12'hE44 : Post_Data = 8'hED; 
	12'hE45 : Post_Data = 8'hED; 
	12'hE46 : Post_Data = 8'hED; 
	12'hE47 : Post_Data = 8'hED; 
	12'hE48 : Post_Data = 8'hED; 
	12'hE49 : Post_Data = 8'hED; 
	12'hE4A : Post_Data = 8'hED; 
	12'hE4B : Post_Data = 8'hED; 
	12'hE4C : Post_Data = 8'hEE; 
	12'hE4D : Post_Data = 8'hEE; 
	12'hE4E : Post_Data = 8'hEE; 
	12'hE4F : Post_Data = 8'hEE; 
	12'hE50 : Post_Data = 8'hEE; 
	12'hE51 : Post_Data = 8'hEE; 
	12'hE52 : Post_Data = 8'hEE; 
	12'hE53 : Post_Data = 8'hEE; 
	12'hE54 : Post_Data = 8'hEE; 
	12'hE55 : Post_Data = 8'hEE; 
	12'hE56 : Post_Data = 8'hEE; 
	12'hE57 : Post_Data = 8'hEE; 
	12'hE58 : Post_Data = 8'hEE; 
	12'hE59 : Post_Data = 8'hEE; 
	12'hE5A : Post_Data = 8'hEE; 
	12'hE5B : Post_Data = 8'hEE; 
	12'hE5C : Post_Data = 8'hEE; 
	12'hE5D : Post_Data = 8'hEE; 
	12'hE5E : Post_Data = 8'hEE; 
	12'hE5F : Post_Data = 8'hEE; 
	12'hE60 : Post_Data = 8'hEE; 
	12'hE61 : Post_Data = 8'hEE; 
	12'hE62 : Post_Data = 8'hEE; 
	12'hE63 : Post_Data = 8'hEF; 
	12'hE64 : Post_Data = 8'hEF; 
	12'hE65 : Post_Data = 8'hEF; 
	12'hE66 : Post_Data = 8'hEF; 
	12'hE67 : Post_Data = 8'hEF; 
	12'hE68 : Post_Data = 8'hEF; 
	12'hE69 : Post_Data = 8'hEF; 
	12'hE6A : Post_Data = 8'hEF; 
	12'hE6B : Post_Data = 8'hEF; 
	12'hE6C : Post_Data = 8'hEF; 
	12'hE6D : Post_Data = 8'hEF; 
	12'hE6E : Post_Data = 8'hEF; 
	12'hE6F : Post_Data = 8'hEF; 
	12'hE70 : Post_Data = 8'hEF; 
	12'hE71 : Post_Data = 8'hEF; 
	12'hE72 : Post_Data = 8'hEF; 
	12'hE73 : Post_Data = 8'hEF; 
	12'hE74 : Post_Data = 8'hEF; 
	12'hE75 : Post_Data = 8'hEF; 
	12'hE76 : Post_Data = 8'hEF; 
	12'hE77 : Post_Data = 8'hEF; 
	12'hE78 : Post_Data = 8'hEF; 
	12'hE79 : Post_Data = 8'hEF; 
	12'hE7A : Post_Data = 8'hF0; 
	12'hE7B : Post_Data = 8'hF0; 
	12'hE7C : Post_Data = 8'hF0; 
	12'hE7D : Post_Data = 8'hF0; 
	12'hE7E : Post_Data = 8'hF0; 
	12'hE7F : Post_Data = 8'hF0; 
	12'hE80 : Post_Data = 8'hF0; 
	12'hE81 : Post_Data = 8'hF0; 
	12'hE82 : Post_Data = 8'hF0; 
	12'hE83 : Post_Data = 8'hF0; 
	12'hE84 : Post_Data = 8'hF0; 
	12'hE85 : Post_Data = 8'hF0; 
	12'hE86 : Post_Data = 8'hF0; 
	12'hE87 : Post_Data = 8'hF0; 
	12'hE88 : Post_Data = 8'hF0; 
	12'hE89 : Post_Data = 8'hF0; 
	12'hE8A : Post_Data = 8'hF0; 
	12'hE8B : Post_Data = 8'hF0; 
	12'hE8C : Post_Data = 8'hF0; 
	12'hE8D : Post_Data = 8'hF0; 
	12'hE8E : Post_Data = 8'hF0; 
	12'hE8F : Post_Data = 8'hF0; 
	12'hE90 : Post_Data = 8'hF0; 
	12'hE91 : Post_Data = 8'hF1; 
	12'hE92 : Post_Data = 8'hF1; 
	12'hE93 : Post_Data = 8'hF1; 
	12'hE94 : Post_Data = 8'hF1; 
	12'hE95 : Post_Data = 8'hF1; 
	12'hE96 : Post_Data = 8'hF1; 
	12'hE97 : Post_Data = 8'hF1; 
	12'hE98 : Post_Data = 8'hF1; 
	12'hE99 : Post_Data = 8'hF1; 
	12'hE9A : Post_Data = 8'hF1; 
	12'hE9B : Post_Data = 8'hF1; 
	12'hE9C : Post_Data = 8'hF1; 
	12'hE9D : Post_Data = 8'hF1; 
	12'hE9E : Post_Data = 8'hF1; 
	12'hE9F : Post_Data = 8'hF1; 
	12'hEA0 : Post_Data = 8'hF1; 
	12'hEA1 : Post_Data = 8'hF1; 
	12'hEA2 : Post_Data = 8'hF1; 
	12'hEA3 : Post_Data = 8'hF1; 
	12'hEA4 : Post_Data = 8'hF1; 
	12'hEA5 : Post_Data = 8'hF1; 
	12'hEA6 : Post_Data = 8'hF1; 
	12'hEA7 : Post_Data = 8'hF1; 
	12'hEA8 : Post_Data = 8'hF2; 
	12'hEA9 : Post_Data = 8'hF2; 
	12'hEAA : Post_Data = 8'hF2; 
	12'hEAB : Post_Data = 8'hF2; 
	12'hEAC : Post_Data = 8'hF2; 
	12'hEAD : Post_Data = 8'hF2; 
	12'hEAE : Post_Data = 8'hF2; 
	12'hEAF : Post_Data = 8'hF2; 
	12'hEB0 : Post_Data = 8'hF2; 
	12'hEB1 : Post_Data = 8'hF2; 
	12'hEB2 : Post_Data = 8'hF2; 
	12'hEB3 : Post_Data = 8'hF2; 
	12'hEB4 : Post_Data = 8'hF2; 
	12'hEB5 : Post_Data = 8'hF2; 
	12'hEB6 : Post_Data = 8'hF2; 
	12'hEB7 : Post_Data = 8'hF2; 
	12'hEB8 : Post_Data = 8'hF2; 
	12'hEB9 : Post_Data = 8'hF2; 
	12'hEBA : Post_Data = 8'hF2; 
	12'hEBB : Post_Data = 8'hF2; 
	12'hEBC : Post_Data = 8'hF2; 
	12'hEBD : Post_Data = 8'hF2; 
	12'hEBE : Post_Data = 8'hF2; 
	12'hEBF : Post_Data = 8'hF2; 
	12'hEC0 : Post_Data = 8'hF3; 
	12'hEC1 : Post_Data = 8'hF3; 
	12'hEC2 : Post_Data = 8'hF3; 
	12'hEC3 : Post_Data = 8'hF3; 
	12'hEC4 : Post_Data = 8'hF3; 
	12'hEC5 : Post_Data = 8'hF3; 
	12'hEC6 : Post_Data = 8'hF3; 
	12'hEC7 : Post_Data = 8'hF3; 
	12'hEC8 : Post_Data = 8'hF3; 
	12'hEC9 : Post_Data = 8'hF3; 
	12'hECA : Post_Data = 8'hF3; 
	12'hECB : Post_Data = 8'hF3; 
	12'hECC : Post_Data = 8'hF3; 
	12'hECD : Post_Data = 8'hF3; 
	12'hECE : Post_Data = 8'hF3; 
	12'hECF : Post_Data = 8'hF3; 
	12'hED0 : Post_Data = 8'hF3; 
	12'hED1 : Post_Data = 8'hF3; 
	12'hED2 : Post_Data = 8'hF3; 
	12'hED3 : Post_Data = 8'hF3; 
	12'hED4 : Post_Data = 8'hF3; 
	12'hED5 : Post_Data = 8'hF3; 
	12'hED6 : Post_Data = 8'hF3; 
	12'hED7 : Post_Data = 8'hF4; 
	12'hED8 : Post_Data = 8'hF4; 
	12'hED9 : Post_Data = 8'hF4; 
	12'hEDA : Post_Data = 8'hF4; 
	12'hEDB : Post_Data = 8'hF4; 
	12'hEDC : Post_Data = 8'hF4; 
	12'hEDD : Post_Data = 8'hF4; 
	12'hEDE : Post_Data = 8'hF4; 
	12'hEDF : Post_Data = 8'hF4; 
	12'hEE0 : Post_Data = 8'hF4; 
	12'hEE1 : Post_Data = 8'hF4; 
	12'hEE2 : Post_Data = 8'hF4; 
	12'hEE3 : Post_Data = 8'hF4; 
	12'hEE4 : Post_Data = 8'hF4; 
	12'hEE5 : Post_Data = 8'hF4; 
	12'hEE6 : Post_Data = 8'hF4; 
	12'hEE7 : Post_Data = 8'hF4; 
	12'hEE8 : Post_Data = 8'hF4; 
	12'hEE9 : Post_Data = 8'hF4; 
	12'hEEA : Post_Data = 8'hF4; 
	12'hEEB : Post_Data = 8'hF4; 
	12'hEEC : Post_Data = 8'hF4; 
	12'hEED : Post_Data = 8'hF4; 
	12'hEEE : Post_Data = 8'hF4; 
	12'hEEF : Post_Data = 8'hF5; 
	12'hEF0 : Post_Data = 8'hF5; 
	12'hEF1 : Post_Data = 8'hF5; 
	12'hEF2 : Post_Data = 8'hF5; 
	12'hEF3 : Post_Data = 8'hF5; 
	12'hEF4 : Post_Data = 8'hF5; 
	12'hEF5 : Post_Data = 8'hF5; 
	12'hEF6 : Post_Data = 8'hF5; 
	12'hEF7 : Post_Data = 8'hF5; 
	12'hEF8 : Post_Data = 8'hF5; 
	12'hEF9 : Post_Data = 8'hF5; 
	12'hEFA : Post_Data = 8'hF5; 
	12'hEFB : Post_Data = 8'hF5; 
	12'hEFC : Post_Data = 8'hF5; 
	12'hEFD : Post_Data = 8'hF5; 
	12'hEFE : Post_Data = 8'hF5; 
	12'hEFF : Post_Data = 8'hF5; 
	12'hF00 : Post_Data = 8'hF5; 
	12'hF01 : Post_Data = 8'hF5; 
	12'hF02 : Post_Data = 8'hF5; 
	12'hF03 : Post_Data = 8'hF5; 
	12'hF04 : Post_Data = 8'hF5; 
	12'hF05 : Post_Data = 8'hF5; 
	12'hF06 : Post_Data = 8'hF6; 
	12'hF07 : Post_Data = 8'hF6; 
	12'hF08 : Post_Data = 8'hF6; 
	12'hF09 : Post_Data = 8'hF6; 
	12'hF0A : Post_Data = 8'hF6; 
	12'hF0B : Post_Data = 8'hF6; 
	12'hF0C : Post_Data = 8'hF6; 
	12'hF0D : Post_Data = 8'hF6; 
	12'hF0E : Post_Data = 8'hF6; 
	12'hF0F : Post_Data = 8'hF6; 
	12'hF10 : Post_Data = 8'hF6; 
	12'hF11 : Post_Data = 8'hF6; 
	12'hF12 : Post_Data = 8'hF6; 
	12'hF13 : Post_Data = 8'hF6; 
	12'hF14 : Post_Data = 8'hF6; 
	12'hF15 : Post_Data = 8'hF6; 
	12'hF16 : Post_Data = 8'hF6; 
	12'hF17 : Post_Data = 8'hF6; 
	12'hF18 : Post_Data = 8'hF6; 
	12'hF19 : Post_Data = 8'hF6; 
	12'hF1A : Post_Data = 8'hF6; 
	12'hF1B : Post_Data = 8'hF6; 
	12'hF1C : Post_Data = 8'hF6; 
	12'hF1D : Post_Data = 8'hF6; 
	12'hF1E : Post_Data = 8'hF7; 
	12'hF1F : Post_Data = 8'hF7; 
	12'hF20 : Post_Data = 8'hF7; 
	12'hF21 : Post_Data = 8'hF7; 
	12'hF22 : Post_Data = 8'hF7; 
	12'hF23 : Post_Data = 8'hF7; 
	12'hF24 : Post_Data = 8'hF7; 
	12'hF25 : Post_Data = 8'hF7; 
	12'hF26 : Post_Data = 8'hF7; 
	12'hF27 : Post_Data = 8'hF7; 
	12'hF28 : Post_Data = 8'hF7; 
	12'hF29 : Post_Data = 8'hF7; 
	12'hF2A : Post_Data = 8'hF7; 
	12'hF2B : Post_Data = 8'hF7; 
	12'hF2C : Post_Data = 8'hF7; 
	12'hF2D : Post_Data = 8'hF7; 
	12'hF2E : Post_Data = 8'hF7; 
	12'hF2F : Post_Data = 8'hF7; 
	12'hF30 : Post_Data = 8'hF7; 
	12'hF31 : Post_Data = 8'hF7; 
	12'hF32 : Post_Data = 8'hF7; 
	12'hF33 : Post_Data = 8'hF7; 
	12'hF34 : Post_Data = 8'hF7; 
	12'hF35 : Post_Data = 8'hF8; 
	12'hF36 : Post_Data = 8'hF8; 
	12'hF37 : Post_Data = 8'hF8; 
	12'hF38 : Post_Data = 8'hF8; 
	12'hF39 : Post_Data = 8'hF8; 
	12'hF3A : Post_Data = 8'hF8; 
	12'hF3B : Post_Data = 8'hF8; 
	12'hF3C : Post_Data = 8'hF8; 
	12'hF3D : Post_Data = 8'hF8; 
	12'hF3E : Post_Data = 8'hF8; 
	12'hF3F : Post_Data = 8'hF8; 
	12'hF40 : Post_Data = 8'hF8; 
	12'hF41 : Post_Data = 8'hF8; 
	12'hF42 : Post_Data = 8'hF8; 
	12'hF43 : Post_Data = 8'hF8; 
	12'hF44 : Post_Data = 8'hF8; 
	12'hF45 : Post_Data = 8'hF8; 
	12'hF46 : Post_Data = 8'hF8; 
	12'hF47 : Post_Data = 8'hF8; 
	12'hF48 : Post_Data = 8'hF8; 
	12'hF49 : Post_Data = 8'hF8; 
	12'hF4A : Post_Data = 8'hF8; 
	12'hF4B : Post_Data = 8'hF8; 
	12'hF4C : Post_Data = 8'hF8; 
	12'hF4D : Post_Data = 8'hF9; 
	12'hF4E : Post_Data = 8'hF9; 
	12'hF4F : Post_Data = 8'hF9; 
	12'hF50 : Post_Data = 8'hF9; 
	12'hF51 : Post_Data = 8'hF9; 
	12'hF52 : Post_Data = 8'hF9; 
	12'hF53 : Post_Data = 8'hF9; 
	12'hF54 : Post_Data = 8'hF9; 
	12'hF55 : Post_Data = 8'hF9; 
	12'hF56 : Post_Data = 8'hF9; 
	12'hF57 : Post_Data = 8'hF9; 
	12'hF58 : Post_Data = 8'hF9; 
	12'hF59 : Post_Data = 8'hF9; 
	12'hF5A : Post_Data = 8'hF9; 
	12'hF5B : Post_Data = 8'hF9; 
	12'hF5C : Post_Data = 8'hF9; 
	12'hF5D : Post_Data = 8'hF9; 
	12'hF5E : Post_Data = 8'hF9; 
	12'hF5F : Post_Data = 8'hF9; 
	12'hF60 : Post_Data = 8'hF9; 
	12'hF61 : Post_Data = 8'hF9; 
	12'hF62 : Post_Data = 8'hF9; 
	12'hF63 : Post_Data = 8'hF9; 
	12'hF64 : Post_Data = 8'hFA; 
	12'hF65 : Post_Data = 8'hFA; 
	12'hF66 : Post_Data = 8'hFA; 
	12'hF67 : Post_Data = 8'hFA; 
	12'hF68 : Post_Data = 8'hFA; 
	12'hF69 : Post_Data = 8'hFA; 
	12'hF6A : Post_Data = 8'hFA; 
	12'hF6B : Post_Data = 8'hFA; 
	12'hF6C : Post_Data = 8'hFA; 
	12'hF6D : Post_Data = 8'hFA; 
	12'hF6E : Post_Data = 8'hFA; 
	12'hF6F : Post_Data = 8'hFA; 
	12'hF70 : Post_Data = 8'hFA; 
	12'hF71 : Post_Data = 8'hFA; 
	12'hF72 : Post_Data = 8'hFA; 
	12'hF73 : Post_Data = 8'hFA; 
	12'hF74 : Post_Data = 8'hFA; 
	12'hF75 : Post_Data = 8'hFA; 
	12'hF76 : Post_Data = 8'hFA; 
	12'hF77 : Post_Data = 8'hFA; 
	12'hF78 : Post_Data = 8'hFA; 
	12'hF79 : Post_Data = 8'hFA; 
	12'hF7A : Post_Data = 8'hFA; 
	12'hF7B : Post_Data = 8'hFA; 
	12'hF7C : Post_Data = 8'hFB; 
	12'hF7D : Post_Data = 8'hFB; 
	12'hF7E : Post_Data = 8'hFB; 
	12'hF7F : Post_Data = 8'hFB; 
	12'hF80 : Post_Data = 8'hFB; 
	12'hF81 : Post_Data = 8'hFB; 
	12'hF82 : Post_Data = 8'hFB; 
	12'hF83 : Post_Data = 8'hFB; 
	12'hF84 : Post_Data = 8'hFB; 
	12'hF85 : Post_Data = 8'hFB; 
	12'hF86 : Post_Data = 8'hFB; 
	12'hF87 : Post_Data = 8'hFB; 
	12'hF88 : Post_Data = 8'hFB; 
	12'hF89 : Post_Data = 8'hFB; 
	12'hF8A : Post_Data = 8'hFB; 
	12'hF8B : Post_Data = 8'hFB; 
	12'hF8C : Post_Data = 8'hFB; 
	12'hF8D : Post_Data = 8'hFB; 
	12'hF8E : Post_Data = 8'hFB; 
	12'hF8F : Post_Data = 8'hFB; 
	12'hF90 : Post_Data = 8'hFB; 
	12'hF91 : Post_Data = 8'hFB; 
	12'hF92 : Post_Data = 8'hFB; 
	12'hF93 : Post_Data = 8'hFB; 
	12'hF94 : Post_Data = 8'hFC; 
	12'hF95 : Post_Data = 8'hFC; 
	12'hF96 : Post_Data = 8'hFC; 
	12'hF97 : Post_Data = 8'hFC; 
	12'hF98 : Post_Data = 8'hFC; 
	12'hF99 : Post_Data = 8'hFC; 
	12'hF9A : Post_Data = 8'hFC; 
	12'hF9B : Post_Data = 8'hFC; 
	12'hF9C : Post_Data = 8'hFC; 
	12'hF9D : Post_Data = 8'hFC; 
	12'hF9E : Post_Data = 8'hFC; 
	12'hF9F : Post_Data = 8'hFC; 
	12'hFA0 : Post_Data = 8'hFC; 
	12'hFA1 : Post_Data = 8'hFC; 
	12'hFA2 : Post_Data = 8'hFC; 
	12'hFA3 : Post_Data = 8'hFC; 
	12'hFA4 : Post_Data = 8'hFC; 
	12'hFA5 : Post_Data = 8'hFC; 
	12'hFA6 : Post_Data = 8'hFC; 
	12'hFA7 : Post_Data = 8'hFC; 
	12'hFA8 : Post_Data = 8'hFC; 
	12'hFA9 : Post_Data = 8'hFC; 
	12'hFAA : Post_Data = 8'hFC; 
	12'hFAB : Post_Data = 8'hFC; 
	12'hFAC : Post_Data = 8'hFD; 
	12'hFAD : Post_Data = 8'hFD; 
	12'hFAE : Post_Data = 8'hFD; 
	12'hFAF : Post_Data = 8'hFD; 
	12'hFB0 : Post_Data = 8'hFD; 
	12'hFB1 : Post_Data = 8'hFD; 
	12'hFB2 : Post_Data = 8'hFD; 
	12'hFB3 : Post_Data = 8'hFD; 
	12'hFB4 : Post_Data = 8'hFD; 
	12'hFB5 : Post_Data = 8'hFD; 
	12'hFB6 : Post_Data = 8'hFD; 
	12'hFB7 : Post_Data = 8'hFD; 
	12'hFB8 : Post_Data = 8'hFD; 
	12'hFB9 : Post_Data = 8'hFD; 
	12'hFBA : Post_Data = 8'hFD; 
	12'hFBB : Post_Data = 8'hFD; 
	12'hFBC : Post_Data = 8'hFD; 
	12'hFBD : Post_Data = 8'hFD; 
	12'hFBE : Post_Data = 8'hFD; 
	12'hFBF : Post_Data = 8'hFD; 
	12'hFC0 : Post_Data = 8'hFD; 
	12'hFC1 : Post_Data = 8'hFD; 
	12'hFC2 : Post_Data = 8'hFD; 
	12'hFC3 : Post_Data = 8'hFD; 
	12'hFC4 : Post_Data = 8'hFE; 
	12'hFC5 : Post_Data = 8'hFE; 
	12'hFC6 : Post_Data = 8'hFE; 
	12'hFC7 : Post_Data = 8'hFE; 
	12'hFC8 : Post_Data = 8'hFE; 
	12'hFC9 : Post_Data = 8'hFE; 
	12'hFCA : Post_Data = 8'hFE; 
	12'hFCB : Post_Data = 8'hFE; 
	12'hFCC : Post_Data = 8'hFE; 
	12'hFCD : Post_Data = 8'hFE; 
	12'hFCE : Post_Data = 8'hFE; 
	12'hFCF : Post_Data = 8'hFE; 
	12'hFD0 : Post_Data = 8'hFE; 
	12'hFD1 : Post_Data = 8'hFE; 
	12'hFD2 : Post_Data = 8'hFE; 
	12'hFD3 : Post_Data = 8'hFE; 
	12'hFD4 : Post_Data = 8'hFE; 
	12'hFD5 : Post_Data = 8'hFE; 
	12'hFD6 : Post_Data = 8'hFE; 
	12'hFD7 : Post_Data = 8'hFE; 
	12'hFD8 : Post_Data = 8'hFE; 
	12'hFD9 : Post_Data = 8'hFE; 
	12'hFDA : Post_Data = 8'hFE; 
	12'hFDB : Post_Data = 8'hFE; 
	12'hFDC : Post_Data = 8'hFF; 
	12'hFDD : Post_Data = 8'hFF; 
	12'hFDE : Post_Data = 8'hFF; 
	12'hFDF : Post_Data = 8'hFF; 
	12'hFE0 : Post_Data = 8'hFF; 
	12'hFE1 : Post_Data = 8'hFF; 
	12'hFE2 : Post_Data = 8'hFF; 
	12'hFE3 : Post_Data = 8'hFF; 
	12'hFE4 : Post_Data = 8'hFF; 
	12'hFE5 : Post_Data = 8'hFF; 
	12'hFE6 : Post_Data = 8'hFF; 
	12'hFE7 : Post_Data = 8'hFF; 
	12'hFE8 : Post_Data = 8'hFF; 
	12'hFE9 : Post_Data = 8'hFF; 
	12'hFEA : Post_Data = 8'hFF; 
	12'hFEB : Post_Data = 8'hFF; 
	12'hFEC : Post_Data = 8'hFF; 
	12'hFED : Post_Data = 8'hFF; 
	12'hFEE : Post_Data = 8'hFF; 
	12'hFEF : Post_Data = 8'hFF; 
	12'hFF0 : Post_Data = 8'hFF; 
	12'hFF1 : Post_Data = 8'hFF; 
	12'hFF2 : Post_Data = 8'hFF; 
	12'hFF3 : Post_Data = 8'hFF; 
	12'hFF4 : Post_Data = 8'hFF; 
	12'hFF5 : Post_Data = 8'hFF; 
	12'hFF6 : Post_Data = 8'hFF; 
	12'hFF7 : Post_Data = 8'hFF; 
	12'hFF8 : Post_Data = 8'hFF; 
	12'hFF9 : Post_Data = 8'hFF; 
	12'hFFA : Post_Data = 8'hFF; 
	12'hFFB : Post_Data = 8'hFF; 
	12'hFFC : Post_Data = 8'hFF; 
	12'hFFD : Post_Data = 8'hFF; 
	12'hFFE : Post_Data = 8'hFF; 
	12'hFFF : Post_Data = 8'hFF; 
	endcase
end

endmodule
